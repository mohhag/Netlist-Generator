
//Verilog file of module FIR


`timescale 1 ns / 1ns

module FIR_net(reset,
clk,
x,
y);
	input reset;
	input clk;
input [0:7]x;
output [0:7]y;
wire
wire_1,
wire_2,
wire_3,
wire_4,
wire_5,
wire_6,
wire_7,
wire_8,
wire_9,
wire_10,
wire_11,
wire_12,
wire_13,
wire_14,
wire_15,
wire_16,
wire_17,
wire_18,
wire_19,
wire_20,
wire_21,
wire_22,
wire_23,
wire_24,
wire_25,
wire_26,
wire_27,
wire_28,
wire_29,
wire_30,
wire_31,
wire_32,
wire_33,
wire_34,
wire_35,
wire_36,
wire_37,
wire_38,
wire_39,
wire_40,
wire_41,
wire_42,
wire_43,
wire_44,
wire_45,
wire_46,
wire_47,
wire_48,
wire_49,
wire_50,
wire_51,
wire_52,
wire_53,
wire_54,
wire_55,
wire_56,
wire_57,
wire_58,
wire_59,
wire_60,
wire_61,
wire_62,
wire_63,
wire_64,
wire_65,
wire_66,
wire_67,
wire_68,
wire_69,
wire_70,
wire_71,
wire_72,
wire_73,
wire_74,
wire_75,
wire_76,
wire_77,
wire_78,
wire_79,
wire_80,
wire_81,
wire_82,
wire_83,
wire_84,
wire_85,
wire_86,
wire_87,
wire_88,
wire_89,
wire_90,
wire_91,
wire_92,
wire_93,
wire_94,
wire_95,
wire_96,
wire_97,
wire_98,
wire_99,
wire_100,
wire_101,
wire_102,
wire_103,
wire_104,
wire_105,
wire_106,
wire_107,
wire_108,
wire_109,
wire_110,
wire_111,
wire_112,
wire_113,
wire_114,
wire_115,
wire_116,
wire_117,
wire_118,
wire_119,
wire_120,
wire_121,
wire_122,
wire_123,
wire_124,
wire_125,
wire_126,
wire_127,
wire_128,
wire_129,
wire_130,
wire_131,
wire_132,
wire_133,
wire_134,
wire_135,
wire_136,
wire_137,
wire_138,
wire_139,
wire_140,
wire_141,
wire_142,
wire_143,
wire_144,
wire_145,
wire_146,
wire_147,
wire_148,
wire_149,
wire_150,
wire_151,
wire_152,
wire_153,
wire_154,
wire_155,
wire_156,
wire_157,
wire_158,
wire_159,
wire_160,
wire_161,
wire_162,
wire_163,
wire_164,
wire_165,
wire_166,
wire_167,
wire_168,
wire_169,
wire_170,
wire_171,
wire_172,
wire_173,
wire_174,
wire_175,
wire_176,
wire_177,
wire_178,
wire_179,
wire_180,
wire_181,
wire_182,
wire_183,
wire_184,
wire_185,
wire_186,
wire_187,
wire_188,
wire_189,
wire_190,
wire_191,
wire_192,
wire_193,
wire_194,
wire_195,
wire_196,
wire_197,
wire_198,
wire_199,
wire_200,
wire_201,
wire_202,
wire_203,
wire_204,
wire_205,
wire_206,
wire_207,
wire_208,
wire_209,
wire_210,
wire_211,
wire_212,
wire_213,
wire_214,
wire_215,
wire_216,
wire_217,
wire_218,
wire_219,
wire_220,
wire_221,
wire_222,
wire_223,
wire_224,
wire_225,
wire_226,
wire_227,
wire_228,
wire_229,
wire_230,
wire_231,
wire_232,
wire_233,
wire_234,
wire_235,
wire_236,
wire_237,
wire_238,
wire_239,
wire_240,
wire_241,
wire_242,
wire_243,
wire_244,
wire_245,
wire_246,
wire_247,
wire_248,
wire_249,
wire_250,
wire_251,
wire_252,
wire_253,
wire_254,
wire_255,
wire_256,
wire_257,
wire_258,
wire_259,
wire_260,
wire_261,
wire_262,
wire_263,
wire_264,
wire_265,
wire_266,
wire_267,
wire_268,
wire_269,
wire_270,
wire_271,
wire_272,
wire_273,
wire_274,
wire_275,
wire_276,
wire_277,
wire_278,
wire_279,
wire_280,
wire_281,
wire_282,
wire_283,
wire_284,
wire_285,
wire_286,
wire_287,
wire_288,
wire_289,
wire_290,
wire_291,
wire_292,
wire_293,
wire_294,
wire_295,
wire_296,
wire_297,
wire_298,
wire_299,
wire_300,
wire_301,
wire_302,
wire_303,
wire_304,
wire_305,
wire_306,
wire_307,
wire_308,
wire_309,
wire_310,
wire_311,
wire_312,
wire_313,
wire_314,
wire_315,
wire_316,
wire_317,
wire_318,
wire_319,
wire_320,
wire_321,
wire_322,
wire_323,
wire_324,
wire_325,
wire_326,
wire_327,
wire_328,
wire_329,
wire_330,
wire_331,
wire_332,
wire_333,
wire_334,
wire_335,
wire_336,
wire_337,
wire_338,
wire_339,
wire_340,
wire_341,
wire_342,
wire_343,
wire_344,
wire_345,
wire_346,
wire_347,
wire_348,
wire_349,
wire_350,
wire_351,
wire_352,
wire_353,
wire_354,
wire_355,
wire_356,
wire_357,
wire_358,
wire_359,
wire_360,
wire_361,
wire_362,
wire_363,
wire_364,
wire_365,
wire_366,
wire_367,
wire_368,
wire_369,
wire_370,
wire_371,
wire_372,
wire_373,
wire_374,
wire_375,
wire_376,
wire_377,
wire_378,
wire_379,
wire_380,
wire_381,
wire_382,
wire_383,
wire_384,
wire_385,
wire_386,
wire_387,
wire_388,
wire_389,
wire_390,
wire_391,
wire_392,
wire_393,
wire_394,
wire_395,
wire_396,
wire_397,
wire_398,
wire_399,
wire_400,
wire_401,
wire_402,
wire_403,
wire_404,
wire_405,
wire_406,
wire_407,
wire_408,
wire_409,
wire_410,
wire_411,
wire_412,
wire_413,
wire_414,
wire_415,
wire_416,
wire_417,
wire_418,
wire_419,
wire_420,
wire_421,
wire_422,
wire_423,
wire_424,
wire_425,
wire_426,
wire_427,
wire_428,
wire_429,
wire_430,
wire_431,
wire_432,
wire_433,
wire_434,
wire_435,
wire_436,
wire_437,
wire_438,
wire_439,
wire_440,
wire_441,
wire_442,
wire_443,
wire_444,
wire_445,
wire_446,
wire_447,
wire_448,
wire_449,
wire_450,
wire_451,
wire_452,
wire_453,
wire_454,
wire_455,
wire_456,
wire_457,
wire_458,
wire_459,
wire_460,
wire_461,
wire_462,
wire_463,
wire_464,
wire_465,
wire_466,
wire_467,
wire_468,
wire_469,
wire_470,
wire_471,
wire_472,
wire_473,
wire_474,
wire_475,
wire_476,
wire_477,
wire_478,
wire_479,
wire_480,
wire_481,
wire_482,
wire_483,
wire_484,
wire_485,
wire_486,
wire_487,
wire_488,
wire_489,
wire_490,
wire_491,
wire_492,
wire_493,
wire_494,
wire_495,
wire_496,
wire_497,
wire_498,
wire_499,
wire_500,
wire_501,
wire_502,
wire_503,
wire_504,
wire_505,
wire_506,
wire_507,
wire_508,
wire_509,
wire_510,
wire_511,
wire_512,
wire_513,
wire_514,
wire_515,
wire_516,
wire_517,
wire_518,
wire_519,
wire_520,
wire_521,
wire_522,
wire_523,
wire_524,
wire_525,
wire_526,
wire_527,
wire_528,
wire_529,
wire_530,
wire_531,
wire_532,
wire_533,
wire_534,
wire_535,
wire_536,
wire_537,
wire_538,
wire_539,
wire_540,
wire_541,
wire_542,
wire_543,
wire_544,
wire_545,
wire_546,
wire_547,
wire_548,
wire_549,
wire_550,
wire_551,
wire_552,
wire_553,
wire_554,
wire_555,
wire_556,
wire_557,
wire_558,
wire_559,
wire_560,
wire_561,
wire_562,
wire_563,
wire_564,
wire_565,
wire_566,
wire_567,
wire_568,
wire_569,
wire_570,
wire_571,
wire_572,
wire_573,
wire_574,
wire_575,
wire_576,
wire_577,
wire_578,
wire_579,
wire_580,
wire_581,
wire_582,
wire_583,
wire_584,
wire_585,
wire_586,
wire_587,
wire_588,
wire_589,
wire_590,
wire_591,
wire_592,
wire_593,
wire_594,
wire_595,
wire_596,
wire_597,
wire_598,
wire_599,
wire_600,
wire_601,
wire_602,
wire_603,
wire_604,
wire_605,
wire_606,
wire_607,
wire_608,
wire_609,
wire_610,
wire_611,
wire_612,
wire_613,
wire_614,
wire_615,
wire_616,
wire_617,
wire_618,
wire_619,
wire_620,
wire_621,
wire_622,
wire_623,
wire_624,
wire_625,
wire_626,
wire_627,
wire_628,
wire_629,
wire_630,
wire_631,
wire_632,
wire_633,
wire_634,
wire_635,
wire_636,
wire_637,
wire_638,
wire_639,
wire_640,
wire_641,
wire_642,
wire_643,
wire_644,
wire_645,
wire_646,
wire_647,
wire_648,
wire_649,
wire_650,
wire_651,
wire_652,
wire_653,
wire_654,
wire_655,
wire_656,
wire_657,
wire_658,
wire_659,
wire_660,
wire_661,
wire_662,
wire_663,
wire_664,
wire_665,
wire_666,
wire_667,
wire_668,
wire_669,
wire_670,
wire_671,
wire_672,
wire_673,
wire_674,
wire_675,
wire_676,
wire_677,
wire_678,
wire_679,
wire_680,
wire_681,
wire_682,
wire_683,
wire_684,
wire_685,
wire_686,
wire_687,
wire_688,
wire_689,
wire_690,
wire_691,
wire_692,
wire_693,
wire_694,
wire_695,
wire_696,
wire_697,
wire_698,
wire_699,
wire_700,
wire_701,
wire_702,
wire_703,
wire_704,
wire_705,
wire_706,
wire_707,
wire_708,
wire_709,
wire_710,
wire_711,
wire_712,
wire_713,
wire_714,
wire_715,
wire_716,
wire_717,
wire_718,
wire_719,
wire_720,
wire_721,
wire_722,
wire_723,
wire_724,
wire_725,
wire_726,
wire_727,
wire_728,
wire_729,
wire_730,
wire_731,
wire_732,
wire_733,
wire_734,
wire_735,
wire_736,
wire_737,
wire_738,
wire_739,
wire_740,
wire_741,
wire_742,
wire_743,
wire_744,
wire_745,
wire_746,
wire_747,
wire_748,
wire_749,
wire_750,
wire_751,
wire_752,
wire_753,
wire_754,
wire_755,
wire_756,
wire_757,
wire_758,
wire_759,
wire_760,
wire_761,
wire_762,
wire_763,
wire_764,
wire_765,
wire_766,
wire_767,
wire_768,
wire_769,
wire_770,
wire_771,
wire_772,
wire_773,
wire_774,
wire_775,
wire_776,
wire_777,
wire_778,
wire_779,
wire_780,
wire_781,
wire_782,
wire_783,
wire_784,
wire_785,
wire_786,
wire_787,
wire_788,
wire_789,
wire_790,
wire_791,
wire_792,
wire_793,
wire_794,
wire_795,
wire_796,
wire_797,
wire_798,
wire_799,
wire_800,
wire_801,
wire_802,
wire_803,
wire_804,
wire_805,
wire_806,
wire_807,
wire_808,
wire_809,
wire_810,
wire_811,
wire_812,
wire_813,
wire_814,
wire_815,
wire_816,
wire_817,
wire_818,
wire_819,
wire_820,
wire_821,
wire_822,
wire_823,
wire_824,
wire_825,
wire_826,
wire_827,
wire_828,
wire_829,
wire_830,
wire_831,
wire_832,
wire_833,
wire_834,
wire_835,
wire_836,
wire_837,
wire_838,
wire_839,
wire_840,
wire_841,
wire_842,
wire_843,
wire_844,
wire_845,
wire_846,
wire_847,
wire_848,
wire_849,
wire_850,
wire_851,
wire_852,
wire_853,
wire_854,
wire_855,
wire_856,
wire_857,
wire_858,
wire_859,
wire_860,
wire_861,
wire_862,
wire_863,
wire_864,
wire_865,
wire_866,
wire_867,
wire_868,
wire_869,
wire_870,
wire_871,
wire_872,
wire_873,
wire_874,
wire_875,
wire_876,
wire_877,
wire_878,
wire_879,
wire_880,
wire_881,
wire_882,
wire_883,
wire_884,
wire_885,
wire_886,
wire_887,
wire_888,
wire_889,
wire_890,
wire_891,
wire_892,
wire_893,
wire_894,
wire_895,
wire_896,
wire_897,
wire_898,
wire_899,
wire_900,
wire_901,
wire_902,
wire_903,
wire_904,
wire_905,
wire_906,
wire_907,
wire_908,
wire_909,
wire_910,
wire_911,
wire_912,
wire_913,
wire_914,
wire_915,
wire_916,
wire_917,
wire_918,
wire_919,
wire_920,
wire_921,
wire_922,
wire_923,
wire_924,
wire_925,
wire_926,
wire_927,
wire_928,
wire_929,
wire_930,
wire_931,
wire_932,
wire_933,
wire_934,
wire_935,
wire_936,
wire_937,
wire_938,
wire_939,
wire_940,
wire_941,
wire_942,
wire_943,
wire_944,
wire_945,
wire_946,
wire_947,
wire_948,
wire_949,
wire_950,
wire_951,
wire_952,
wire_953,
wire_954,
wire_955,
wire_956,
wire_957,
wire_958,
wire_959,
wire_960,
wire_961,
wire_962,
wire_963,
wire_964,
wire_965,
wire_966,
wire_967,
wire_968,
wire_969,
wire_970,
wire_971,
wire_972,
wire_973,
wire_974,
wire_975,
wire_976,
wire_977,
wire_978,
wire_979,
wire_980,
wire_981,
wire_982,
wire_983,
wire_984,
wire_985,
wire_986,
wire_987,
wire_988,
wire_989,
wire_990,
wire_991,
wire_992,
wire_993,
wire_994,
wire_995,
wire_996,
wire_997,
wire_998,
wire_999,
wire_1000,
wire_1001,
wire_1002,
wire_1003,
wire_1004,
wire_1005,
wire_1006,
wire_1007,
wire_1008,
wire_1009,
wire_1010,
wire_1011,
wire_1012,
wire_1013,
wire_1014,
wire_1015,
wire_1016,
wire_1017,
wire_1018,
wire_1019,
wire_1020,
wire_1021,
wire_1022,
wire_1023,
wire_1024,
wire_1025,
wire_1026,
wire_1027,
wire_1028,
wire_1029,
wire_1030,
wire_1031,
wire_1032,
wire_1033,
wire_1034,
wire_1035,
wire_1036,
wire_1037,
wire_1038,
wire_1039,
wire_1040,
wire_1041,
wire_1042,
wire_1043,
wire_1044,
wire_1045,
wire_1046,
wire_1047,
wire_1048,
wire_1049,
wire_1050,
wire_1051,
wire_1052,
wire_1053,
wire_1054,
wire_1055,
wire_1056,
wire_1057,
wire_1058,
wire_1059,
wire_1060,
wire_1061,
wire_1062,
wire_1063,
wire_1064,
wire_1065,
wire_1066,
wire_1067,
wire_1068,
wire_1069,
wire_1070,
wire_1071,
wire_1072,
wire_1073,
wire_1074,
wire_1075,
wire_1076,
wire_1077,
wire_42_0,
wire_42_1,
wire_43_0,
wire_43_1,
wire_43_2,
wire_44_0,
wire_44_1,
wire_44_2,
wire_45_0,
wire_45_1,
wire_45_2,
wire_46_0,
wire_46_1,
wire_46_2,
wire_47_0,
wire_47_1,
wire_47_2,
wire_48_0,
wire_48_1,
wire_48_2,
wire_90_0,
wire_90_1,
wire_91_0,
wire_91_1,
wire_92_0,
wire_92_1,
wire_93_0,
wire_93_1,
wire_94_0,
wire_94_1,
wire_95_0,
wire_95_1,
wire_96_0,
wire_96_1,
wire_96_2,
wire_123_0,
wire_123_1,
wire_124_0,
wire_124_1,
wire_124_2,
wire_125_0,
wire_125_1,
wire_125_2,
wire_126_0,
wire_126_1,
wire_126_2,
wire_127_0,
wire_127_1,
wire_127_2,
wire_128_0,
wire_128_1,
wire_128_2,
wire_129_0,
wire_129_1,
wire_129_2,
wire_155_0,
wire_155_1,
wire_156_0,
wire_156_1,
wire_157_0,
wire_157_1,
wire_158_0,
wire_158_1,
wire_159_0,
wire_159_1,
wire_160_0,
wire_160_1,
wire_161_0,
wire_161_1,
wire_161_2,
wire_163_0,
wire_163_1,
wire_163_2,
wire_163_3,
wire_163_4,
wire_163_5,
wire_163_6,
wire_193_0,
wire_193_1,
wire_194_0,
wire_194_1,
wire_195_0,
wire_195_1,
wire_196_0,
wire_196_1,
wire_197_0,
wire_197_1,
wire_198_0,
wire_198_1,
wire_200_0,
wire_200_1,
wire_200_2,
wire_200_3,
wire_200_4,
wire_200_5,
wire_241_0,
wire_241_1,
wire_241_2,
wire_242_0,
wire_242_1,
wire_242_2,
wire_243_0,
wire_243_1,
wire_243_2,
wire_244_0,
wire_244_1,
wire_244_2,
wire_245_0,
wire_245_1,
wire_245_2,
wire_246_0,
wire_246_1,
wire_246_2,
wire_247_0,
wire_247_1,
wire_249_0,
wire_249_1,
wire_249_2,
wire_249_3,
wire_249_4,
wire_249_5,
wire_249_6,
wire_249_7,
wire_290_0,
wire_290_1,
wire_290_2,
wire_291_0,
wire_291_1,
wire_291_2,
wire_291_3,
wire_292_0,
wire_292_1,
wire_292_2,
wire_292_3,
wire_293_0,
wire_293_1,
wire_293_2,
wire_293_3,
wire_294_0,
wire_294_1,
wire_294_2,
wire_294_3,
wire_295_0,
wire_295_1,
wire_295_2,
wire_295_3,
wire_296_0,
wire_296_1,
wire_298_0,
wire_298_1,
wire_298_2,
wire_298_3,
wire_298_4,
wire_298_5,
wire_339_0,
wire_339_1,
wire_339_2,
wire_340_0,
wire_340_1,
wire_340_2,
wire_340_3,
wire_341_0,
wire_341_1,
wire_341_2,
wire_341_3,
wire_342_0,
wire_342_1,
wire_342_2,
wire_342_3,
wire_343_0,
wire_343_1,
wire_343_2,
wire_343_3,
wire_344_0,
wire_344_1,
wire_344_2,
wire_344_3,
wire_345_0,
wire_345_1,
wire_345_2,
wire_345_3,
wire_493_0,
wire_493_1,
wire_493_2,
wire_493_3,
wire_493_4,
wire_493_5,
wire_493_6,
wire_493_7,
wire_493_8,
wire_493_9,
wire_493_10,
wire_493_11,
wire_493_12,
wire_493_13,
wire_493_14,
wire_493_15,
wire_383_0,
wire_383_1,
wire_383_2,
wire_383_3,
wire_383_4,
wire_383_5,
wire_383_6,
wire_383_7,
wire_383_8,
wire_383_9,
wire_383_10,
wire_383_11,
wire_383_12,
wire_383_13,
wire_383_14,
wire_680_0,
wire_680_1,
wire_703_0,
wire_703_1,
wire_703_2,
wire_704_0,
wire_704_1,
wire_704_2,
wire_699_0,
wire_699_1,
wire_699_2,
wire_694_0,
wire_694_1,
wire_694_2,
wire_689_0,
wire_689_1,
wire_689_2,
wire_690_0,
wire_690_1,
wire_695_0,
wire_695_1,
wire_700_0,
wire_700_1,
wire_705_0,
wire_705_1,
wire_679_0,
wire_679_1,
wire_698_0,
wire_698_1,
wire_698_2,
wire_693_0,
wire_693_1,
wire_693_2,
wire_688_0,
wire_688_1,
wire_688_2,
wire_763_0,
wire_763_1,
wire_763_2,
wire_768_0,
wire_768_1,
wire_768_2,
wire_773_0,
wire_773_1,
wire_773_2,
wire_778_0,
wire_778_1,
wire_778_2,
wire_754_0,
wire_754_1,
wire_777_0,
wire_777_1,
wire_777_2,
wire_786_0,
wire_786_1,
wire_786_2,
wire_790_0,
wire_790_1,
wire_794_0,
wire_794_1,
wire_798_0,
wire_798_1,
wire_802_0,
wire_802_1,
wire_801_0,
wire_801_1,
wire_801_2,
wire_752_0,
wire_752_1,
wire_787_0,
wire_787_1,
wire_787_2,
wire_791_0,
wire_791_1,
wire_791_2,
wire_795_0,
wire_795_1,
wire_795_2,
wire_799_0,
wire_799_1,
wire_799_2,
wire_803_0,
wire_803_1,
wire_803_2,
wire_751_0,
wire_751_1,
wire_764_0,
wire_764_1,
wire_769_0,
wire_769_1,
wire_774_0,
wire_774_1,
wire_779_0,
wire_779_1,
wire_753_0,
wire_753_1,
wire_797_0,
wire_797_1,
wire_797_2,
wire_793_0,
wire_793_1,
wire_793_2,
wire_789_0,
wire_789_1,
wire_789_2,
wire_785_0,
wire_785_1,
wire_785_2,
wire_772_0,
wire_772_1,
wire_772_2,
wire_767_0,
wire_767_1,
wire_767_2,
wire_762_0,
wire_762_1,
wire_762_2,
wire_859_0,
wire_859_1,
wire_859_2,
wire_863_0,
wire_863_1,
wire_867_0,
wire_867_1,
wire_871_0,
wire_871_1,
wire_875_0,
wire_875_1,
wire_874_0,
wire_874_1,
wire_874_2,
wire_851_0,
wire_851_1,
wire_870_0,
wire_870_1,
wire_870_2,
wire_866_0,
wire_866_1,
wire_866_2,
wire_862_0,
wire_862_1,
wire_862_2,
wire_858_0,
wire_858_1,
wire_858_2,
wire_932_0,
wire_932_1,
wire_932_2,
wire_937_0,
wire_937_1,
wire_937_2,
wire_942_0,
wire_942_1,
wire_942_2,
wire_947_0,
wire_947_1,
wire_947_2,
wire_923_0,
wire_923_1,
wire_946_0,
wire_946_1,
wire_946_2,
wire_954_0,
wire_954_1,
wire_954_2,
wire_957_0,
wire_957_1,
wire_957_2,
wire_960_0,
wire_960_1,
wire_960_2,
wire_963_0,
wire_963_1,
wire_963_2,
wire_966_0,
wire_966_1,
wire_966_2,
wire_965_0,
wire_965_1,
wire_965_2,
wire_921_0,
wire_921_1,
wire_933_0,
wire_933_1,
wire_938_0,
wire_938_1,
wire_943_0,
wire_943_1,
wire_948_0,
wire_948_1,
wire_922_0,
wire_922_1,
wire_962_0,
wire_962_1,
wire_962_2,
wire_959_0,
wire_959_1,
wire_959_2,
wire_956_0,
wire_956_1,
wire_956_2,
wire_953_0,
wire_953_1,
wire_953_2,
wire_941_0,
wire_941_1,
wire_941_2,
wire_936_0,
wire_936_1,
wire_936_2,
wire_931_0,
wire_931_1,
wire_931_2,
wire_380_0,
wire_380_1,
wire_403_0,
wire_403_1,
wire_400_0,
wire_400_1,
wire_397_0,
wire_397_1,
wire_394_0,
wire_394_1,
wire_391_0,
wire_391_1,
wire_388_0,
wire_388_1,
wire_385_0,
wire_385_1,
wire_1027_0,
wire_1027_1,
wire_1027_2,
wire_1025_0,
wire_1025_1,
wire_1025_2,
wire_1023_0,
wire_1023_1,
wire_1023_2,
wire_1021_0,
wire_1021_1,
wire_1021_2,
wire_1019_0,
wire_1019_1,
wire_1019_2,
wire_1017_0,
wire_1017_1,
wire_1017_2,
wire_348_0,
wire_348_1,
wire_376_0,
wire_376_1,
wire_372_0,
wire_372_1,
wire_368_0,
wire_368_1,
wire_364_0,
wire_364_1,
wire_360_0,
wire_360_1,
wire_356_0,
wire_356_1,
wire_352_0,
wire_352_1,
wire_1059_0,
wire_1059_1,
wire_1059_2,
wire_1057_0,
wire_1057_1,
wire_1057_2,
wire_1055_0,
wire_1055_1,
wire_1055_2,
wire_1053_0,
wire_1053_1,
wire_1053_2,
wire_1051_0,
wire_1051_1,
wire_1051_2,
wire_1049_0,
wire_1049_1,
wire_1049_2,
wire_556_0,
wire_556_1,
wire_556_2,
wire_556_3,
wire_556_4,
wire_556_5,
wire_556_6,
wire_556_7,
wire_556_8,
wire_556_9,
wire_556_10,
wire_556_11,
wire_556_12,
wire_556_13,
wire_556_14,
wire_556_15,
wire_556_16,
wire_556_17,
wire_556_18,
wire_556_19,
wire_556_20,
wire_556_21,
wire_556_22,
wire_556_23,
wire_556_24,
wire_556_25,
wire_556_26,
wire_556_27,
wire_556_28,
wire_556_29,
wire_556_30,
wire_556_31,
wire_556_32,
wire_556_33,
wire_556_34,
wire_556_35,
wire_556_36,
wire_556_37,
wire_556_38,
wire_556_39,
wire_556_40,
wire_556_41,
wire_556_42,
wire_556_43,
wire_556_44,
wire_556_45,
wire_556_46,
wire_556_47,
wire_556_48,
wire_556_49,
wire_556_50,
wire_556_51,
wire_556_52,
wire_556_53,
wire_556_54,
wire_556_55,
wire_556_56,
wire_556_57,
wire_556_58,
wire_556_59,
wire_556_60,
wire_556_61,
wire_556_62,
wire_556_63,
wire_556_64,
wire_556_65,
wire_556_66,
wire_556_67,
wire_556_68,
wire_556_69,
wire_556_70,
wire_556_71,
wire_556_72,
wire_556_73,
wire_556_74,
wire_556_75,
wire_556_76,
wire_556_77,
wire_556_78,
wire_556_79,
wire_556_80,
wire_556_81,
wire_556_82,
wire_556_83,
wire_556_84,
wire_556_85,
wire_556_86,
wire_324_0,
wire_324_1,
wire_326_0,
wire_326_1,
wire_328_0,
wire_328_1,
wire_330_0,
wire_330_1,
wire_332_0,
wire_332_1,
wire_334_0,
wire_334_1,
wire_336_0,
wire_336_1,
wire_338_0,
wire_338_1,
reset_net_0,
clk_net_0;

pin #(10) pin_0 ({reset, clk, x[0], x[1], x[2], x[3], x[4], x[5], x[6], x[7]}, {reset_net_0, clk_net_0, x_0, x_1, x_2, x_3, x_4, x_5, x_6, x_7});

pout #(8) pout_0 ({y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7}, {y[0], y[1], y[2], y[3], y[4], y[5], y[6], y[7]});

fanout_n #(2, 0, 0) FANOUT_1 (wire_42, {wire_42_0, wire_42_1});
fanout_n #(3, 0, 0) FANOUT_2 (wire_43, {wire_43_0, wire_43_1, wire_43_2});
fanout_n #(3, 0, 0) FANOUT_3 (wire_44, {wire_44_0, wire_44_1, wire_44_2});
fanout_n #(3, 0, 0) FANOUT_4 (wire_45, {wire_45_0, wire_45_1, wire_45_2});
fanout_n #(3, 0, 0) FANOUT_5 (wire_46, {wire_46_0, wire_46_1, wire_46_2});
fanout_n #(3, 0, 0) FANOUT_6 (wire_47, {wire_47_0, wire_47_1, wire_47_2});
fanout_n #(3, 0, 0) FANOUT_7 (wire_48, {wire_48_0, wire_48_1, wire_48_2});
fanout_n #(2, 0, 0) FANOUT_8 (wire_90, {wire_90_0, wire_90_1});
fanout_n #(2, 0, 0) FANOUT_9 (wire_91, {wire_91_0, wire_91_1});
fanout_n #(2, 0, 0) FANOUT_10 (wire_92, {wire_92_0, wire_92_1});
fanout_n #(2, 0, 0) FANOUT_11 (wire_93, {wire_93_0, wire_93_1});
fanout_n #(2, 0, 0) FANOUT_12 (wire_94, {wire_94_0, wire_94_1});
fanout_n #(2, 0, 0) FANOUT_13 (wire_95, {wire_95_0, wire_95_1});
fanout_n #(3, 0, 0) FANOUT_14 (wire_96, {wire_96_0, wire_96_1, wire_96_2});
fanout_n #(2, 0, 0) FANOUT_15 (wire_123, {wire_123_0, wire_123_1});
fanout_n #(3, 0, 0) FANOUT_16 (wire_124, {wire_124_0, wire_124_1, wire_124_2});
fanout_n #(3, 0, 0) FANOUT_17 (wire_125, {wire_125_0, wire_125_1, wire_125_2});
fanout_n #(3, 0, 0) FANOUT_18 (wire_126, {wire_126_0, wire_126_1, wire_126_2});
fanout_n #(3, 0, 0) FANOUT_19 (wire_127, {wire_127_0, wire_127_1, wire_127_2});
fanout_n #(3, 0, 0) FANOUT_20 (wire_128, {wire_128_0, wire_128_1, wire_128_2});
fanout_n #(3, 0, 0) FANOUT_21 (wire_129, {wire_129_0, wire_129_1, wire_129_2});
fanout_n #(2, 0, 0) FANOUT_22 (wire_155, {wire_155_0, wire_155_1});
fanout_n #(2, 0, 0) FANOUT_23 (wire_156, {wire_156_0, wire_156_1});
fanout_n #(2, 0, 0) FANOUT_24 (wire_157, {wire_157_0, wire_157_1});
fanout_n #(2, 0, 0) FANOUT_25 (wire_158, {wire_158_0, wire_158_1});
fanout_n #(2, 0, 0) FANOUT_26 (wire_159, {wire_159_0, wire_159_1});
fanout_n #(2, 0, 0) FANOUT_27 (wire_160, {wire_160_0, wire_160_1});
fanout_n #(3, 0, 0) FANOUT_28 (wire_161, {wire_161_0, wire_161_1, wire_161_2});
fanout_n #(7, 0, 0) FANOUT_29 (wire_163, {wire_163_0, wire_163_1, wire_163_2, wire_163_3, wire_163_4, wire_163_5, wire_163_6});
fanout_n #(2, 0, 0) FANOUT_30 (wire_193, {wire_193_0, wire_193_1});
fanout_n #(2, 0, 0) FANOUT_31 (wire_194, {wire_194_0, wire_194_1});
fanout_n #(2, 0, 0) FANOUT_32 (wire_195, {wire_195_0, wire_195_1});
fanout_n #(2, 0, 0) FANOUT_33 (wire_196, {wire_196_0, wire_196_1});
fanout_n #(2, 0, 0) FANOUT_34 (wire_197, {wire_197_0, wire_197_1});
fanout_n #(2, 0, 0) FANOUT_35 (wire_198, {wire_198_0, wire_198_1});
fanout_n #(6, 0, 0) FANOUT_36 (wire_200, {wire_200_0, wire_200_1, wire_200_2, wire_200_3, wire_200_4, wire_200_5});
fanout_n #(3, 0, 0) FANOUT_37 (wire_241, {wire_241_0, wire_241_1, wire_241_2});
fanout_n #(3, 0, 0) FANOUT_38 (wire_242, {wire_242_0, wire_242_1, wire_242_2});
fanout_n #(3, 0, 0) FANOUT_39 (wire_243, {wire_243_0, wire_243_1, wire_243_2});
fanout_n #(3, 0, 0) FANOUT_40 (wire_244, {wire_244_0, wire_244_1, wire_244_2});
fanout_n #(3, 0, 0) FANOUT_41 (wire_245, {wire_245_0, wire_245_1, wire_245_2});
fanout_n #(3, 0, 0) FANOUT_42 (wire_246, {wire_246_0, wire_246_1, wire_246_2});
fanout_n #(2, 0, 0) FANOUT_43 (wire_247, {wire_247_0, wire_247_1});
fanout_n #(8, 0, 0) FANOUT_44 (wire_249, {wire_249_0, wire_249_1, wire_249_2, wire_249_3, wire_249_4, wire_249_5, wire_249_6, wire_249_7});
fanout_n #(3, 0, 0) FANOUT_45 (wire_290, {wire_290_0, wire_290_1, wire_290_2});
fanout_n #(4, 0, 0) FANOUT_46 (wire_291, {wire_291_0, wire_291_1, wire_291_2, wire_291_3});
fanout_n #(4, 0, 0) FANOUT_47 (wire_292, {wire_292_0, wire_292_1, wire_292_2, wire_292_3});
fanout_n #(4, 0, 0) FANOUT_48 (wire_293, {wire_293_0, wire_293_1, wire_293_2, wire_293_3});
fanout_n #(4, 0, 0) FANOUT_49 (wire_294, {wire_294_0, wire_294_1, wire_294_2, wire_294_3});
fanout_n #(4, 0, 0) FANOUT_50 (wire_295, {wire_295_0, wire_295_1, wire_295_2, wire_295_3});
fanout_n #(2, 0, 0) FANOUT_51 (wire_296, {wire_296_0, wire_296_1});
fanout_n #(6, 0, 0) FANOUT_52 (wire_298, {wire_298_0, wire_298_1, wire_298_2, wire_298_3, wire_298_4, wire_298_5});
fanout_n #(3, 0, 0) FANOUT_53 (wire_339, {wire_339_0, wire_339_1, wire_339_2});
fanout_n #(4, 0, 0) FANOUT_54 (wire_340, {wire_340_0, wire_340_1, wire_340_2, wire_340_3});
fanout_n #(4, 0, 0) FANOUT_55 (wire_341, {wire_341_0, wire_341_1, wire_341_2, wire_341_3});
fanout_n #(4, 0, 0) FANOUT_56 (wire_342, {wire_342_0, wire_342_1, wire_342_2, wire_342_3});
fanout_n #(4, 0, 0) FANOUT_57 (wire_343, {wire_343_0, wire_343_1, wire_343_2, wire_343_3});
fanout_n #(4, 0, 0) FANOUT_58 (wire_344, {wire_344_0, wire_344_1, wire_344_2, wire_344_3});
fanout_n #(4, 0, 0) FANOUT_59 (wire_345, {wire_345_0, wire_345_1, wire_345_2, wire_345_3});
fanout_n #(16, 0, 0) FANOUT_60 (wire_493, {wire_493_0, wire_493_1, wire_493_2, wire_493_3, wire_493_4, wire_493_5, wire_493_6, wire_493_7, wire_493_8, wire_493_9, wire_493_10, wire_493_11, wire_493_12, wire_493_13, wire_493_14, wire_493_15});
fanout_n #(15, 0, 0) FANOUT_61 (wire_383, {wire_383_0, wire_383_1, wire_383_2, wire_383_3, wire_383_4, wire_383_5, wire_383_6, wire_383_7, wire_383_8, wire_383_9, wire_383_10, wire_383_11, wire_383_12, wire_383_13, wire_383_14});
fanout_n #(2, 0, 0) FANOUT_62 (wire_680, {wire_680_0, wire_680_1});
fanout_n #(3, 0, 0) FANOUT_63 (wire_703, {wire_703_0, wire_703_1, wire_703_2});
fanout_n #(3, 0, 0) FANOUT_64 (wire_704, {wire_704_0, wire_704_1, wire_704_2});
fanout_n #(3, 0, 0) FANOUT_65 (wire_699, {wire_699_0, wire_699_1, wire_699_2});
fanout_n #(3, 0, 0) FANOUT_66 (wire_694, {wire_694_0, wire_694_1, wire_694_2});
fanout_n #(3, 0, 0) FANOUT_67 (wire_689, {wire_689_0, wire_689_1, wire_689_2});
fanout_n #(2, 0, 0) FANOUT_68 (wire_690, {wire_690_0, wire_690_1});
fanout_n #(2, 0, 0) FANOUT_69 (wire_695, {wire_695_0, wire_695_1});
fanout_n #(2, 0, 0) FANOUT_70 (wire_700, {wire_700_0, wire_700_1});
fanout_n #(2, 0, 0) FANOUT_71 (wire_705, {wire_705_0, wire_705_1});
fanout_n #(2, 0, 0) FANOUT_72 (wire_679, {wire_679_0, wire_679_1});
fanout_n #(3, 0, 0) FANOUT_73 (wire_698, {wire_698_0, wire_698_1, wire_698_2});
fanout_n #(3, 0, 0) FANOUT_74 (wire_693, {wire_693_0, wire_693_1, wire_693_2});
fanout_n #(3, 0, 0) FANOUT_75 (wire_688, {wire_688_0, wire_688_1, wire_688_2});
fanout_n #(3, 0, 0) FANOUT_76 (wire_763, {wire_763_0, wire_763_1, wire_763_2});
fanout_n #(3, 0, 0) FANOUT_77 (wire_768, {wire_768_0, wire_768_1, wire_768_2});
fanout_n #(3, 0, 0) FANOUT_78 (wire_773, {wire_773_0, wire_773_1, wire_773_2});
fanout_n #(3, 0, 0) FANOUT_79 (wire_778, {wire_778_0, wire_778_1, wire_778_2});
fanout_n #(2, 0, 0) FANOUT_80 (wire_754, {wire_754_0, wire_754_1});
fanout_n #(3, 0, 0) FANOUT_81 (wire_777, {wire_777_0, wire_777_1, wire_777_2});
fanout_n #(3, 0, 0) FANOUT_82 (wire_786, {wire_786_0, wire_786_1, wire_786_2});
fanout_n #(2, 0, 0) FANOUT_83 (wire_790, {wire_790_0, wire_790_1});
fanout_n #(2, 0, 0) FANOUT_84 (wire_794, {wire_794_0, wire_794_1});
fanout_n #(2, 0, 0) FANOUT_85 (wire_798, {wire_798_0, wire_798_1});
fanout_n #(2, 0, 0) FANOUT_86 (wire_802, {wire_802_0, wire_802_1});
fanout_n #(3, 0, 0) FANOUT_87 (wire_801, {wire_801_0, wire_801_1, wire_801_2});
fanout_n #(2, 0, 0) FANOUT_88 (wire_752, {wire_752_0, wire_752_1});
fanout_n #(3, 0, 0) FANOUT_89 (wire_787, {wire_787_0, wire_787_1, wire_787_2});
fanout_n #(3, 0, 0) FANOUT_90 (wire_791, {wire_791_0, wire_791_1, wire_791_2});
fanout_n #(3, 0, 0) FANOUT_91 (wire_795, {wire_795_0, wire_795_1, wire_795_2});
fanout_n #(3, 0, 0) FANOUT_92 (wire_799, {wire_799_0, wire_799_1, wire_799_2});
fanout_n #(3, 0, 0) FANOUT_93 (wire_803, {wire_803_0, wire_803_1, wire_803_2});
fanout_n #(2, 0, 0) FANOUT_94 (wire_751, {wire_751_0, wire_751_1});
fanout_n #(2, 0, 0) FANOUT_95 (wire_764, {wire_764_0, wire_764_1});
fanout_n #(2, 0, 0) FANOUT_96 (wire_769, {wire_769_0, wire_769_1});
fanout_n #(2, 0, 0) FANOUT_97 (wire_774, {wire_774_0, wire_774_1});
fanout_n #(2, 0, 0) FANOUT_98 (wire_779, {wire_779_0, wire_779_1});
fanout_n #(2, 0, 0) FANOUT_99 (wire_753, {wire_753_0, wire_753_1});
fanout_n #(3, 0, 0) FANOUT_100 (wire_797, {wire_797_0, wire_797_1, wire_797_2});
fanout_n #(3, 0, 0) FANOUT_101 (wire_793, {wire_793_0, wire_793_1, wire_793_2});
fanout_n #(3, 0, 0) FANOUT_102 (wire_789, {wire_789_0, wire_789_1, wire_789_2});
fanout_n #(3, 0, 0) FANOUT_103 (wire_785, {wire_785_0, wire_785_1, wire_785_2});
fanout_n #(3, 0, 0) FANOUT_104 (wire_772, {wire_772_0, wire_772_1, wire_772_2});
fanout_n #(3, 0, 0) FANOUT_105 (wire_767, {wire_767_0, wire_767_1, wire_767_2});
fanout_n #(3, 0, 0) FANOUT_106 (wire_762, {wire_762_0, wire_762_1, wire_762_2});
fanout_n #(3, 0, 0) FANOUT_107 (wire_859, {wire_859_0, wire_859_1, wire_859_2});
fanout_n #(2, 0, 0) FANOUT_108 (wire_863, {wire_863_0, wire_863_1});
fanout_n #(2, 0, 0) FANOUT_109 (wire_867, {wire_867_0, wire_867_1});
fanout_n #(2, 0, 0) FANOUT_110 (wire_871, {wire_871_0, wire_871_1});
fanout_n #(2, 0, 0) FANOUT_111 (wire_875, {wire_875_0, wire_875_1});
fanout_n #(3, 0, 0) FANOUT_112 (wire_874, {wire_874_0, wire_874_1, wire_874_2});
fanout_n #(2, 0, 0) FANOUT_113 (wire_851, {wire_851_0, wire_851_1});
fanout_n #(3, 0, 0) FANOUT_114 (wire_870, {wire_870_0, wire_870_1, wire_870_2});
fanout_n #(3, 0, 0) FANOUT_115 (wire_866, {wire_866_0, wire_866_1, wire_866_2});
fanout_n #(3, 0, 0) FANOUT_116 (wire_862, {wire_862_0, wire_862_1, wire_862_2});
fanout_n #(3, 0, 0) FANOUT_117 (wire_858, {wire_858_0, wire_858_1, wire_858_2});
fanout_n #(3, 0, 0) FANOUT_118 (wire_932, {wire_932_0, wire_932_1, wire_932_2});
fanout_n #(3, 0, 0) FANOUT_119 (wire_937, {wire_937_0, wire_937_1, wire_937_2});
fanout_n #(3, 0, 0) FANOUT_120 (wire_942, {wire_942_0, wire_942_1, wire_942_2});
fanout_n #(3, 0, 0) FANOUT_121 (wire_947, {wire_947_0, wire_947_1, wire_947_2});
fanout_n #(2, 0, 0) FANOUT_122 (wire_923, {wire_923_0, wire_923_1});
fanout_n #(3, 0, 0) FANOUT_123 (wire_946, {wire_946_0, wire_946_1, wire_946_2});
fanout_n #(3, 0, 0) FANOUT_124 (wire_954, {wire_954_0, wire_954_1, wire_954_2});
fanout_n #(3, 0, 0) FANOUT_125 (wire_957, {wire_957_0, wire_957_1, wire_957_2});
fanout_n #(3, 0, 0) FANOUT_126 (wire_960, {wire_960_0, wire_960_1, wire_960_2});
fanout_n #(3, 0, 0) FANOUT_127 (wire_963, {wire_963_0, wire_963_1, wire_963_2});
fanout_n #(3, 0, 0) FANOUT_128 (wire_966, {wire_966_0, wire_966_1, wire_966_2});
fanout_n #(3, 0, 0) FANOUT_129 (wire_965, {wire_965_0, wire_965_1, wire_965_2});
fanout_n #(2, 0, 0) FANOUT_130 (wire_921, {wire_921_0, wire_921_1});
fanout_n #(2, 0, 0) FANOUT_131 (wire_933, {wire_933_0, wire_933_1});
fanout_n #(2, 0, 0) FANOUT_132 (wire_938, {wire_938_0, wire_938_1});
fanout_n #(2, 0, 0) FANOUT_133 (wire_943, {wire_943_0, wire_943_1});
fanout_n #(2, 0, 0) FANOUT_134 (wire_948, {wire_948_0, wire_948_1});
fanout_n #(2, 0, 0) FANOUT_135 (wire_922, {wire_922_0, wire_922_1});
fanout_n #(3, 0, 0) FANOUT_136 (wire_962, {wire_962_0, wire_962_1, wire_962_2});
fanout_n #(3, 0, 0) FANOUT_137 (wire_959, {wire_959_0, wire_959_1, wire_959_2});
fanout_n #(3, 0, 0) FANOUT_138 (wire_956, {wire_956_0, wire_956_1, wire_956_2});
fanout_n #(3, 0, 0) FANOUT_139 (wire_953, {wire_953_0, wire_953_1, wire_953_2});
fanout_n #(3, 0, 0) FANOUT_140 (wire_941, {wire_941_0, wire_941_1, wire_941_2});
fanout_n #(3, 0, 0) FANOUT_141 (wire_936, {wire_936_0, wire_936_1, wire_936_2});
fanout_n #(3, 0, 0) FANOUT_142 (wire_931, {wire_931_0, wire_931_1, wire_931_2});
fanout_n #(2, 0, 0) FANOUT_143 (wire_380, {wire_380_0, wire_380_1});
fanout_n #(2, 0, 0) FANOUT_144 (wire_403, {wire_403_0, wire_403_1});
fanout_n #(2, 0, 0) FANOUT_145 (wire_400, {wire_400_0, wire_400_1});
fanout_n #(2, 0, 0) FANOUT_146 (wire_397, {wire_397_0, wire_397_1});
fanout_n #(2, 0, 0) FANOUT_147 (wire_394, {wire_394_0, wire_394_1});
fanout_n #(2, 0, 0) FANOUT_148 (wire_391, {wire_391_0, wire_391_1});
fanout_n #(2, 0, 0) FANOUT_149 (wire_388, {wire_388_0, wire_388_1});
fanout_n #(2, 0, 0) FANOUT_150 (wire_385, {wire_385_0, wire_385_1});
fanout_n #(3, 0, 0) FANOUT_151 (wire_1027, {wire_1027_0, wire_1027_1, wire_1027_2});
fanout_n #(3, 0, 0) FANOUT_152 (wire_1025, {wire_1025_0, wire_1025_1, wire_1025_2});
fanout_n #(3, 0, 0) FANOUT_153 (wire_1023, {wire_1023_0, wire_1023_1, wire_1023_2});
fanout_n #(3, 0, 0) FANOUT_154 (wire_1021, {wire_1021_0, wire_1021_1, wire_1021_2});
fanout_n #(3, 0, 0) FANOUT_155 (wire_1019, {wire_1019_0, wire_1019_1, wire_1019_2});
fanout_n #(3, 0, 0) FANOUT_156 (wire_1017, {wire_1017_0, wire_1017_1, wire_1017_2});
fanout_n #(2, 0, 0) FANOUT_157 (wire_348, {wire_348_0, wire_348_1});
fanout_n #(2, 0, 0) FANOUT_158 (wire_376, {wire_376_0, wire_376_1});
fanout_n #(2, 0, 0) FANOUT_159 (wire_372, {wire_372_0, wire_372_1});
fanout_n #(2, 0, 0) FANOUT_160 (wire_368, {wire_368_0, wire_368_1});
fanout_n #(2, 0, 0) FANOUT_161 (wire_364, {wire_364_0, wire_364_1});
fanout_n #(2, 0, 0) FANOUT_162 (wire_360, {wire_360_0, wire_360_1});
fanout_n #(2, 0, 0) FANOUT_163 (wire_356, {wire_356_0, wire_356_1});
fanout_n #(2, 0, 0) FANOUT_164 (wire_352, {wire_352_0, wire_352_1});
fanout_n #(3, 0, 0) FANOUT_165 (wire_1059, {wire_1059_0, wire_1059_1, wire_1059_2});
fanout_n #(3, 0, 0) FANOUT_166 (wire_1057, {wire_1057_0, wire_1057_1, wire_1057_2});
fanout_n #(3, 0, 0) FANOUT_167 (wire_1055, {wire_1055_0, wire_1055_1, wire_1055_2});
fanout_n #(3, 0, 0) FANOUT_168 (wire_1053, {wire_1053_0, wire_1053_1, wire_1053_2});
fanout_n #(3, 0, 0) FANOUT_169 (wire_1051, {wire_1051_0, wire_1051_1, wire_1051_2});
fanout_n #(3, 0, 0) FANOUT_170 (wire_1049, {wire_1049_0, wire_1049_1, wire_1049_2});
fanout_n #(87, 0, 0) FANOUT_171 (wire_556, {wire_556_0, wire_556_1, wire_556_2, wire_556_3, wire_556_4, wire_556_5, wire_556_6, wire_556_7, wire_556_8, wire_556_9, wire_556_10, wire_556_11, wire_556_12, wire_556_13, wire_556_14, wire_556_15, wire_556_16, wire_556_17, wire_556_18, wire_556_19, wire_556_20, wire_556_21, wire_556_22, wire_556_23, wire_556_24, wire_556_25, wire_556_26, wire_556_27, wire_556_28, wire_556_29, wire_556_30, wire_556_31, wire_556_32, wire_556_33, wire_556_34, wire_556_35, wire_556_36, wire_556_37, wire_556_38, wire_556_39, wire_556_40, wire_556_41, wire_556_42, wire_556_43, wire_556_44, wire_556_45, wire_556_46, wire_556_47, wire_556_48, wire_556_49, wire_556_50, wire_556_51, wire_556_52, wire_556_53, wire_556_54, wire_556_55, wire_556_56, wire_556_57, wire_556_58, wire_556_59, wire_556_60, wire_556_61, wire_556_62, wire_556_63, wire_556_64, wire_556_65, wire_556_66, wire_556_67, wire_556_68, wire_556_69, wire_556_70, wire_556_71, wire_556_72, wire_556_73, wire_556_74, wire_556_75, wire_556_76, wire_556_77, wire_556_78, wire_556_79, wire_556_80, wire_556_81, wire_556_82, wire_556_83, wire_556_84, wire_556_85, wire_556_86});
fanout_n #(2, 0, 0) FANOUT_172 (wire_324, {wire_324_0, wire_324_1});
fanout_n #(2, 0, 0) FANOUT_173 (wire_326, {wire_326_0, wire_326_1});
fanout_n #(2, 0, 0) FANOUT_174 (wire_328, {wire_328_0, wire_328_1});
fanout_n #(2, 0, 0) FANOUT_175 (wire_330, {wire_330_0, wire_330_1});
fanout_n #(2, 0, 0) FANOUT_176 (wire_332, {wire_332_0, wire_332_1});
fanout_n #(2, 0, 0) FANOUT_177 (wire_334, {wire_334_0, wire_334_1});
fanout_n #(2, 0, 0) FANOUT_178 (wire_336, {wire_336_0, wire_336_1});
fanout_n #(2, 0, 0) FANOUT_179 (wire_338, {wire_338_0, wire_338_1});


and_n #(2, 0, 0) AND_1 (wire_1, {wire_2, wire_3});
and_n #(2, 0, 0) AND_2 (wire_4, {wire_5, wire_6});
and_n #(2, 0, 0) AND_3 (wire_7, {wire_8, wire_9});
and_n #(2, 0, 0) AND_4 (wire_10, {wire_11, wire_12});
and_n #(2, 0, 0) AND_5 (wire_13, {wire_14, wire_15});
and_n #(2, 0, 0) AND_6 (wire_16, {wire_17, wire_18});
and_n #(2, 0, 0) AND_7 (wire_19, {wire_20, wire_21});
and_n #(2, 0, 0) AND_8 (wire_22, {wire_23, wire_24});
and_n #(2, 0, 0) AND_9 (wire_25, {wire_26, wire_27});
and_n #(2, 0, 0) AND_10 (wire_28, {wire_29, wire_27});
and_n #(2, 0, 0) AND_11 (wire_30, {wire_31, wire_27});
and_n #(2, 0, 0) AND_12 (wire_32, {wire_33, wire_27});
and_n #(2, 0, 0) AND_13 (wire_34, {wire_35, wire_27});
and_n #(2, 0, 0) AND_14 (wire_36, {wire_37, wire_27});
and_n #(2, 0, 0) AND_15 (wire_38, {wire_39, wire_27});
and_n #(2, 0, 0) AND_16 (wire_40, {wire_41, wire_27});
or_n #(2, 0, 0) OR_1 (wire_42, {wire_25, wire_1});
notg #(0, 0) NOT_1 (wire_3, wire_27);
or_n #(2, 0, 0) OR_2 (wire_43, {wire_28, wire_4});
notg #(0, 0) NOT_2 (wire_6, wire_27);
or_n #(2, 0, 0) OR_3 (wire_44, {wire_30, wire_7});
notg #(0, 0) NOT_3 (wire_9, wire_27);
or_n #(2, 0, 0) OR_4 (wire_45, {wire_32, wire_10});
notg #(0, 0) NOT_4 (wire_12, wire_27);
or_n #(2, 0, 0) OR_5 (wire_46, {wire_34, wire_13});
notg #(0, 0) NOT_5 (wire_15, wire_27);
or_n #(2, 0, 0) OR_6 (wire_47, {wire_36, wire_16});
notg #(0, 0) NOT_6 (wire_18, wire_27);
or_n #(2, 0, 0) OR_7 (wire_48, {wire_38, wire_19});
notg #(0, 0) NOT_7 (wire_21, wire_27);
or_n #(2, 0, 0) OR_8 (wire_49, {wire_40, wire_22});
notg #(0, 0) NOT_8 (wire_24, wire_27);
and_n #(2, 0, 0) AND_17 (wire_50, {wire_51, wire_52});
and_n #(2, 0, 0) AND_18 (wire_53, {wire_54, wire_55});
and_n #(2, 0, 0) AND_19 (wire_56, {wire_57, wire_58});
and_n #(2, 0, 0) AND_20 (wire_59, {wire_60, wire_61});
and_n #(2, 0, 0) AND_21 (wire_62, {wire_63, wire_64});
and_n #(2, 0, 0) AND_22 (wire_65, {wire_66, wire_67});
and_n #(2, 0, 0) AND_23 (wire_68, {wire_69, wire_70});
and_n #(2, 0, 0) AND_24 (wire_71, {wire_72, wire_73});
and_n #(2, 0, 0) AND_25 (wire_74, {wire_75, wire_27});
and_n #(2, 0, 0) AND_26 (wire_76, {wire_77, wire_27});
and_n #(2, 0, 0) AND_27 (wire_78, {wire_79, wire_27});
and_n #(2, 0, 0) AND_28 (wire_80, {wire_81, wire_27});
and_n #(2, 0, 0) AND_29 (wire_82, {wire_83, wire_27});
and_n #(2, 0, 0) AND_30 (wire_84, {wire_85, wire_27});
and_n #(2, 0, 0) AND_31 (wire_86, {wire_87, wire_27});
and_n #(2, 0, 0) AND_32 (wire_88, {wire_89, wire_27});
or_n #(2, 0, 0) OR_9 (wire_90, {wire_74, wire_50});
notg #(0, 0) NOT_9 (wire_52, wire_27);
or_n #(2, 0, 0) OR_10 (wire_91, {wire_76, wire_53});
notg #(0, 0) NOT_10 (wire_55, wire_27);
or_n #(2, 0, 0) OR_11 (wire_92, {wire_78, wire_56});
notg #(0, 0) NOT_11 (wire_58, wire_27);
or_n #(2, 0, 0) OR_12 (wire_93, {wire_80, wire_59});
notg #(0, 0) NOT_12 (wire_61, wire_27);
or_n #(2, 0, 0) OR_13 (wire_94, {wire_82, wire_62});
notg #(0, 0) NOT_13 (wire_64, wire_27);
or_n #(2, 0, 0) OR_14 (wire_95, {wire_84, wire_65});
notg #(0, 0) NOT_14 (wire_67, wire_27);
or_n #(2, 0, 0) OR_15 (wire_96, {wire_86, wire_68});
notg #(0, 0) NOT_15 (wire_70, wire_27);
or_n #(2, 0, 0) OR_16 (wire_97, {wire_88, wire_71});
notg #(0, 0) NOT_16 (wire_73, wire_27);
and_n #(2, 0, 0) AND_33 (wire_98, {wire_2, wire_99});
and_n #(2, 0, 0) AND_34 (wire_100, {wire_5, wire_101});
and_n #(2, 0, 0) AND_35 (wire_102, {wire_8, wire_103});
and_n #(2, 0, 0) AND_36 (wire_104, {wire_11, wire_105});
and_n #(2, 0, 0) AND_37 (wire_106, {wire_14, wire_107});
and_n #(2, 0, 0) AND_38 (wire_108, {wire_17, wire_109});
and_n #(2, 0, 0) AND_39 (wire_110, {wire_20, wire_111});
and_n #(2, 0, 0) AND_40 (wire_112, {wire_23, wire_113});
and_n #(2, 0, 0) AND_41 (wire_114, {wire_26, wire_115});
and_n #(2, 0, 0) AND_42 (wire_116, {wire_29, wire_115});
and_n #(2, 0, 0) AND_43 (wire_117, {wire_31, wire_115});
and_n #(2, 0, 0) AND_44 (wire_118, {wire_33, wire_115});
and_n #(2, 0, 0) AND_45 (wire_119, {wire_35, wire_115});
and_n #(2, 0, 0) AND_46 (wire_120, {wire_37, wire_115});
and_n #(2, 0, 0) AND_47 (wire_121, {wire_39, wire_115});
and_n #(2, 0, 0) AND_48 (wire_122, {wire_41, wire_115});
or_n #(2, 0, 0) OR_17 (wire_123, {wire_114, wire_98});
notg #(0, 0) NOT_17 (wire_99, wire_115);
or_n #(2, 0, 0) OR_18 (wire_124, {wire_116, wire_100});
notg #(0, 0) NOT_18 (wire_101, wire_115);
or_n #(2, 0, 0) OR_19 (wire_125, {wire_117, wire_102});
notg #(0, 0) NOT_19 (wire_103, wire_115);
or_n #(2, 0, 0) OR_20 (wire_126, {wire_118, wire_104});
notg #(0, 0) NOT_20 (wire_105, wire_115);
or_n #(2, 0, 0) OR_21 (wire_127, {wire_119, wire_106});
notg #(0, 0) NOT_21 (wire_107, wire_115);
or_n #(2, 0, 0) OR_22 (wire_128, {wire_120, wire_108});
notg #(0, 0) NOT_22 (wire_109, wire_115);
or_n #(2, 0, 0) OR_23 (wire_129, {wire_121, wire_110});
notg #(0, 0) NOT_23 (wire_111, wire_115);
or_n #(2, 0, 0) OR_24 (wire_130, {wire_122, wire_112});
notg #(0, 0) NOT_24 (wire_113, wire_115);
and_n #(2, 0, 0) AND_49 (wire_131, {wire_51, wire_132});
and_n #(2, 0, 0) AND_50 (wire_133, {wire_54, wire_134});
and_n #(2, 0, 0) AND_51 (wire_135, {wire_57, wire_136});
and_n #(2, 0, 0) AND_52 (wire_137, {wire_60, wire_138});
and_n #(2, 0, 0) AND_53 (wire_139, {wire_63, wire_140});
and_n #(2, 0, 0) AND_54 (wire_141, {wire_66, wire_142});
and_n #(2, 0, 0) AND_55 (wire_143, {wire_69, wire_144});
and_n #(2, 0, 0) AND_56 (wire_145, {wire_72, wire_146});
and_n #(2, 0, 0) AND_57 (wire_147, {wire_75, wire_115});
and_n #(2, 0, 0) AND_58 (wire_148, {wire_77, wire_115});
and_n #(2, 0, 0) AND_59 (wire_149, {wire_79, wire_115});
and_n #(2, 0, 0) AND_60 (wire_150, {wire_81, wire_115});
and_n #(2, 0, 0) AND_61 (wire_151, {wire_83, wire_115});
and_n #(2, 0, 0) AND_62 (wire_152, {wire_85, wire_115});
and_n #(2, 0, 0) AND_63 (wire_153, {wire_87, wire_115});
and_n #(2, 0, 0) AND_64 (wire_154, {wire_89, wire_115});
or_n #(2, 0, 0) OR_25 (wire_155, {wire_147, wire_131});
notg #(0, 0) NOT_25 (wire_132, wire_115);
or_n #(2, 0, 0) OR_26 (wire_156, {wire_148, wire_133});
notg #(0, 0) NOT_26 (wire_134, wire_115);
or_n #(2, 0, 0) OR_27 (wire_157, {wire_149, wire_135});
notg #(0, 0) NOT_27 (wire_136, wire_115);
or_n #(2, 0, 0) OR_28 (wire_158, {wire_150, wire_137});
notg #(0, 0) NOT_28 (wire_138, wire_115);
or_n #(2, 0, 0) OR_29 (wire_159, {wire_151, wire_139});
notg #(0, 0) NOT_29 (wire_140, wire_115);
or_n #(2, 0, 0) OR_30 (wire_160, {wire_152, wire_141});
notg #(0, 0) NOT_30 (wire_142, wire_115);
or_n #(2, 0, 0) OR_31 (wire_161, {wire_153, wire_143});
notg #(0, 0) NOT_31 (wire_144, wire_115);
or_n #(2, 0, 0) OR_32 (wire_162, {wire_154, wire_145});
notg #(0, 0) NOT_32 (wire_146, wire_115);
notg #(0, 0) NOT_33 (wire_163, wire_164);
and_n #(2, 0, 0) AND_65 (wire_165, {wire_75, wire_166});
and_n #(2, 0, 0) AND_66 (wire_167, {wire_77, wire_168});
and_n #(2, 0, 0) AND_67 (wire_169, {wire_79, wire_170});
and_n #(2, 0, 0) AND_68 (wire_171, {wire_81, wire_172});
and_n #(2, 0, 0) AND_69 (wire_173, {wire_83, wire_174});
and_n #(2, 0, 0) AND_70 (wire_175, {wire_85, wire_176});
and_n #(2, 0, 0) AND_71 (wire_177, {wire_87, wire_178});
and_n #(2, 0, 0) AND_72 (wire_179, {wire_180, wire_164});
and_n #(2, 0, 0) AND_73 (wire_181, {wire_182, wire_164});
and_n #(2, 0, 0) AND_74 (wire_183, {wire_184, wire_164});
and_n #(2, 0, 0) AND_75 (wire_185, {wire_186, wire_164});
and_n #(2, 0, 0) AND_76 (wire_187, {wire_188, wire_164});
and_n #(2, 0, 0) AND_77 (wire_189, {wire_190, wire_164});
and_n #(2, 0, 0) AND_78 (wire_191, {wire_192, wire_164});
or_n #(2, 0, 0) OR_33 (wire_193, {wire_179, wire_165});
notg #(0, 0) NOT_34 (wire_166, wire_164);
or_n #(2, 0, 0) OR_34 (wire_194, {wire_181, wire_167});
notg #(0, 0) NOT_35 (wire_168, wire_164);
or_n #(2, 0, 0) OR_35 (wire_195, {wire_183, wire_169});
notg #(0, 0) NOT_36 (wire_170, wire_164);
or_n #(2, 0, 0) OR_36 (wire_196, {wire_185, wire_171});
notg #(0, 0) NOT_37 (wire_172, wire_164);
or_n #(2, 0, 0) OR_37 (wire_197, {wire_187, wire_173});
notg #(0, 0) NOT_38 (wire_174, wire_164);
or_n #(2, 0, 0) OR_38 (wire_198, {wire_189, wire_175});
notg #(0, 0) NOT_39 (wire_176, wire_164);
or_n #(2, 0, 0) OR_39 (wire_199, {wire_191, wire_177});
notg #(0, 0) NOT_40 (wire_178, wire_164);
notg #(0, 0) NOT_41 (wire_200, wire_164);
and_n #(2, 0, 0) AND_79 (wire_201, {wire_202, wire_203});
and_n #(2, 0, 0) AND_80 (wire_204, {wire_205, wire_206});
and_n #(2, 0, 0) AND_81 (wire_207, {wire_208, wire_209});
and_n #(2, 0, 0) AND_82 (wire_210, {wire_211, wire_212});
and_n #(2, 0, 0) AND_83 (wire_213, {wire_214, wire_215});
and_n #(2, 0, 0) AND_84 (wire_216, {wire_217, wire_218});
and_n #(2, 0, 0) AND_85 (wire_219, {wire_220, wire_221});
and_n #(2, 0, 0) AND_86 (wire_222, {wire_223, wire_224});
and_n #(2, 0, 0) AND_87 (wire_225, {wire_226, wire_164});
and_n #(2, 0, 0) AND_88 (wire_227, {wire_228, wire_164});
and_n #(2, 0, 0) AND_89 (wire_229, {wire_230, wire_164});
and_n #(2, 0, 0) AND_90 (wire_231, {wire_232, wire_164});
and_n #(2, 0, 0) AND_91 (wire_233, {wire_234, wire_164});
and_n #(2, 0, 0) AND_92 (wire_235, {wire_236, wire_164});
and_n #(2, 0, 0) AND_93 (wire_237, {wire_238, wire_164});
and_n #(2, 0, 0) AND_94 (wire_239, {wire_240, wire_164});
or_n #(2, 0, 0) OR_40 (wire_241, {wire_225, wire_201});
notg #(0, 0) NOT_42 (wire_203, wire_164);
or_n #(2, 0, 0) OR_41 (wire_242, {wire_227, wire_204});
notg #(0, 0) NOT_43 (wire_206, wire_164);
or_n #(2, 0, 0) OR_42 (wire_243, {wire_229, wire_207});
notg #(0, 0) NOT_44 (wire_209, wire_164);
or_n #(2, 0, 0) OR_43 (wire_244, {wire_231, wire_210});
notg #(0, 0) NOT_45 (wire_212, wire_164);
or_n #(2, 0, 0) OR_44 (wire_245, {wire_233, wire_213});
notg #(0, 0) NOT_46 (wire_215, wire_164);
or_n #(2, 0, 0) OR_45 (wire_246, {wire_235, wire_216});
notg #(0, 0) NOT_47 (wire_218, wire_164);
or_n #(2, 0, 0) OR_46 (wire_247, {wire_237, wire_219});
notg #(0, 0) NOT_48 (wire_221, wire_164);
or_n #(2, 0, 0) OR_47 (wire_248, {wire_239, wire_222});
notg #(0, 0) NOT_49 (wire_224, wire_164);
notg #(0, 0) NOT_50 (wire_249, wire_164);
and_n #(2, 0, 0) AND_95 (wire_250, {wire_251, wire_252});
and_n #(2, 0, 0) AND_96 (wire_253, {wire_254, wire_255});
and_n #(2, 0, 0) AND_97 (wire_256, {wire_257, wire_258});
and_n #(2, 0, 0) AND_98 (wire_259, {wire_260, wire_261});
and_n #(2, 0, 0) AND_99 (wire_262, {wire_263, wire_264});
and_n #(2, 0, 0) AND_100 (wire_265, {wire_266, wire_267});
and_n #(2, 0, 0) AND_101 (wire_268, {wire_269, wire_270});
and_n #(2, 0, 0) AND_102 (wire_271, {wire_272, wire_273});
and_n #(2, 0, 0) AND_103 (wire_274, {wire_275, wire_164});
and_n #(2, 0, 0) AND_104 (wire_276, {wire_277, wire_164});
and_n #(2, 0, 0) AND_105 (wire_278, {wire_279, wire_164});
and_n #(2, 0, 0) AND_106 (wire_280, {wire_281, wire_164});
and_n #(2, 0, 0) AND_107 (wire_282, {wire_283, wire_164});
and_n #(2, 0, 0) AND_108 (wire_284, {wire_285, wire_164});
and_n #(2, 0, 0) AND_109 (wire_286, {wire_287, wire_164});
and_n #(2, 0, 0) AND_110 (wire_288, {wire_289, wire_164});
or_n #(2, 0, 0) OR_48 (wire_290, {wire_274, wire_250});
notg #(0, 0) NOT_51 (wire_252, wire_164);
or_n #(2, 0, 0) OR_49 (wire_291, {wire_276, wire_253});
notg #(0, 0) NOT_52 (wire_255, wire_164);
or_n #(2, 0, 0) OR_50 (wire_292, {wire_278, wire_256});
notg #(0, 0) NOT_53 (wire_258, wire_164);
or_n #(2, 0, 0) OR_51 (wire_293, {wire_280, wire_259});
notg #(0, 0) NOT_54 (wire_261, wire_164);
or_n #(2, 0, 0) OR_52 (wire_294, {wire_282, wire_262});
notg #(0, 0) NOT_55 (wire_264, wire_164);
or_n #(2, 0, 0) OR_53 (wire_295, {wire_284, wire_265});
notg #(0, 0) NOT_56 (wire_267, wire_164);
or_n #(2, 0, 0) OR_54 (wire_296, {wire_286, wire_268});
notg #(0, 0) NOT_57 (wire_270, wire_164);
or_n #(2, 0, 0) OR_55 (wire_297, {wire_288, wire_271});
notg #(0, 0) NOT_58 (wire_273, wire_164);
notg #(0, 0) NOT_59 (wire_298, wire_164);
and_n #(2, 0, 0) AND_111 (wire_299, {wire_300, wire_301});
and_n #(2, 0, 0) AND_112 (wire_302, {wire_303, wire_304});
and_n #(2, 0, 0) AND_113 (wire_305, {wire_306, wire_307});
and_n #(2, 0, 0) AND_114 (wire_308, {wire_309, wire_310});
and_n #(2, 0, 0) AND_115 (wire_311, {wire_312, wire_313});
and_n #(2, 0, 0) AND_116 (wire_314, {wire_315, wire_316});
and_n #(2, 0, 0) AND_117 (wire_317, {wire_318, wire_319});
and_n #(2, 0, 0) AND_118 (wire_320, {wire_321, wire_322});
and_n #(2, 0, 0) AND_119 (wire_323, {wire_324_0, wire_164});
and_n #(2, 0, 0) AND_120 (wire_325, {wire_326_0, wire_164});
and_n #(2, 0, 0) AND_121 (wire_327, {wire_328_0, wire_164});
and_n #(2, 0, 0) AND_122 (wire_329, {wire_330_0, wire_164});
and_n #(2, 0, 0) AND_123 (wire_331, {wire_332_0, wire_164});
and_n #(2, 0, 0) AND_124 (wire_333, {wire_334_0, wire_164});
and_n #(2, 0, 0) AND_125 (wire_335, {wire_336_0, wire_164});
and_n #(2, 0, 0) AND_126 (wire_337, {wire_338_0, wire_164});
or_n #(2, 0, 0) OR_56 (wire_339, {wire_323, wire_299});
notg #(0, 0) NOT_60 (wire_301, wire_164);
or_n #(2, 0, 0) OR_57 (wire_340, {wire_325, wire_302});
notg #(0, 0) NOT_61 (wire_304, wire_164);
or_n #(2, 0, 0) OR_58 (wire_341, {wire_327, wire_305});
notg #(0, 0) NOT_62 (wire_307, wire_164);
or_n #(2, 0, 0) OR_59 (wire_342, {wire_329, wire_308});
notg #(0, 0) NOT_63 (wire_310, wire_164);
or_n #(2, 0, 0) OR_60 (wire_343, {wire_331, wire_311});
notg #(0, 0) NOT_64 (wire_313, wire_164);
or_n #(2, 0, 0) OR_61 (wire_344, {wire_333, wire_314});
notg #(0, 0) NOT_65 (wire_316, wire_164);
or_n #(2, 0, 0) OR_62 (wire_345, {wire_335, wire_317});
notg #(0, 0) NOT_66 (wire_319, wire_164);
or_n #(2, 0, 0) OR_63 (wire_346, {wire_337, wire_320});
notg #(0, 0) NOT_67 (wire_322, wire_164);
and_n #(2, 0, 0) AND_127 (wire_347, {wire_348_0, wire_349});
and_n #(2, 0, 0) AND_128 (wire_350, {wire_348_1, wire_27});
and_n #(2, 0, 0) AND_129 (wire_351, {wire_352_0, wire_353});
and_n #(2, 0, 0) AND_130 (wire_354, {wire_352_1, wire_27});
and_n #(2, 0, 0) AND_131 (wire_355, {wire_356_0, wire_357});
and_n #(2, 0, 0) AND_132 (wire_358, {wire_356_1, wire_27});
and_n #(2, 0, 0) AND_133 (wire_359, {wire_360_0, wire_361});
and_n #(2, 0, 0) AND_134 (wire_362, {wire_360_1, wire_27});
and_n #(2, 0, 0) AND_135 (wire_363, {wire_364_0, wire_365});
and_n #(2, 0, 0) AND_136 (wire_366, {wire_364_1, wire_27});
and_n #(2, 0, 0) AND_137 (wire_367, {wire_368_0, wire_369});
and_n #(2, 0, 0) AND_138 (wire_370, {wire_368_1, wire_27});
and_n #(2, 0, 0) AND_139 (wire_371, {wire_372_0, wire_373});
and_n #(2, 0, 0) AND_140 (wire_374, {wire_372_1, wire_27});
and_n #(2, 0, 0) AND_141 (wire_375, {wire_376_0, wire_377});
and_n #(2, 0, 0) AND_142 (wire_378, {wire_376_1, wire_27});
and_n #(2, 0, 0) AND_143 (wire_379, {wire_380_0, wire_381});
and_n #(2, 0, 0) AND_144 (wire_382, {wire_380_1, wire_383_0});
and_n #(2, 0, 0) AND_145 (wire_384, {wire_385_0, wire_381});
and_n #(2, 0, 0) AND_146 (wire_386, {wire_385_1, wire_383_1});
and_n #(2, 0, 0) AND_147 (wire_387, {wire_388_0, wire_381});
and_n #(2, 0, 0) AND_148 (wire_389, {wire_388_1, wire_383_2});
and_n #(2, 0, 0) AND_149 (wire_390, {wire_391_0, wire_381});
and_n #(2, 0, 0) AND_150 (wire_392, {wire_391_1, wire_383_3});
and_n #(2, 0, 0) AND_151 (wire_393, {wire_394_0, wire_381});
and_n #(2, 0, 0) AND_152 (wire_395, {wire_394_1, wire_383_4});
and_n #(2, 0, 0) AND_153 (wire_396, {wire_397_0, wire_381});
and_n #(2, 0, 0) AND_154 (wire_398, {wire_397_1, wire_383_5});
and_n #(2, 0, 0) AND_155 (wire_399, {wire_400_0, wire_381});
and_n #(2, 0, 0) AND_156 (wire_401, {wire_400_1, wire_383_6});
and_n #(2, 0, 0) AND_157 (wire_402, {wire_403_0, wire_381});
and_n #(2, 0, 0) AND_158 (wire_404, {wire_403_1, wire_383_7});
bufg #(0, 0) BUF_1 (wire_405, 1'b0);
or_n #(2, 0, 0) OR_64 (wire_460, {wire_350, wire_461});
notg #(0, 0) NOT_68 (wire_462, wire_27);
and_n #(2, 0, 0) AND_159 (wire_461, {wire_462, wire_339_0});
or_n #(2, 0, 0) OR_65 (wire_463, {wire_354, wire_464});
notg #(0, 0) NOT_69 (wire_465, wire_27);
and_n #(2, 0, 0) AND_160 (wire_464, {wire_465, wire_466});
or_n #(2, 0, 0) OR_66 (wire_467, {wire_358, wire_468});
notg #(0, 0) NOT_70 (wire_469, wire_27);
and_n #(2, 0, 0) AND_161 (wire_468, {wire_469, wire_470});
or_n #(2, 0, 0) OR_67 (wire_471, {wire_362, wire_472});
notg #(0, 0) NOT_71 (wire_473, wire_27);
and_n #(2, 0, 0) AND_162 (wire_472, {wire_473, wire_474});
or_n #(2, 0, 0) OR_68 (wire_475, {wire_366, wire_476});
notg #(0, 0) NOT_72 (wire_477, wire_27);
and_n #(2, 0, 0) AND_163 (wire_476, {wire_477, wire_478});
or_n #(2, 0, 0) OR_69 (wire_479, {wire_370, wire_480});
notg #(0, 0) NOT_73 (wire_481, wire_27);
and_n #(2, 0, 0) AND_164 (wire_480, {wire_481, wire_482});
or_n #(2, 0, 0) OR_70 (wire_483, {wire_374, wire_484});
notg #(0, 0) NOT_74 (wire_485, wire_27);
and_n #(2, 0, 0) AND_165 (wire_484, {wire_485, wire_486});
or_n #(2, 0, 0) OR_71 (wire_487, {wire_378, wire_488});
notg #(0, 0) NOT_75 (wire_489, wire_27);
and_n #(2, 0, 0) AND_166 (wire_488, {wire_489, wire_490});
or_n #(2, 0, 0) OR_72 (wire_491, {wire_492, wire_347});
and_n #(2, 0, 0) AND_167 (wire_492, {wire_493_0, wire_494});
notg #(0, 0) NOT_76 (wire_349, wire_493_1);
or_n #(2, 0, 0) OR_73 (wire_495, {wire_496, wire_351});
and_n #(2, 0, 0) AND_168 (wire_496, {wire_493_2, wire_497});
notg #(0, 0) NOT_77 (wire_353, wire_493_3);
or_n #(2, 0, 0) OR_74 (wire_498, {wire_499, wire_355});
and_n #(2, 0, 0) AND_169 (wire_499, {wire_493_4, wire_500});
notg #(0, 0) NOT_78 (wire_357, wire_493_5);
or_n #(2, 0, 0) OR_75 (wire_501, {wire_502, wire_359});
and_n #(2, 0, 0) AND_170 (wire_502, {wire_493_6, wire_503});
notg #(0, 0) NOT_79 (wire_361, wire_493_7);
or_n #(2, 0, 0) OR_76 (wire_504, {wire_505, wire_363});
and_n #(2, 0, 0) AND_171 (wire_505, {wire_493_8, wire_506});
notg #(0, 0) NOT_80 (wire_365, wire_493_9);
or_n #(2, 0, 0) OR_77 (wire_507, {wire_508, wire_367});
and_n #(2, 0, 0) AND_172 (wire_508, {wire_493_10, wire_509});
notg #(0, 0) NOT_81 (wire_369, wire_493_11);
or_n #(2, 0, 0) OR_78 (wire_510, {wire_511, wire_371});
and_n #(2, 0, 0) AND_173 (wire_511, {wire_493_12, wire_512});
notg #(0, 0) NOT_82 (wire_373, wire_493_13);
or_n #(2, 0, 0) OR_79 (wire_513, {wire_514, wire_375});
and_n #(2, 0, 0) AND_174 (wire_514, {wire_493_14, wire_515});
notg #(0, 0) NOT_83 (wire_377, wire_493_15);
nor_n #(2, 0, 0) NOR_1 (wire_493, {wire_457, wire_115});
or_n #(2, 0, 0) OR_80 (wire_516, {wire_386, wire_517});
notg #(0, 0) NOT_84 (wire_518, wire_383_8);
and_n #(2, 0, 0) AND_175 (wire_517, {wire_518, wire_519});
or_n #(2, 0, 0) OR_81 (wire_520, {wire_389, wire_521});
notg #(0, 0) NOT_85 (wire_522, wire_383_9);
and_n #(2, 0, 0) AND_176 (wire_521, {wire_522, wire_523});
or_n #(2, 0, 0) OR_82 (wire_524, {wire_392, wire_525});
notg #(0, 0) NOT_86 (wire_526, wire_383_10);
and_n #(2, 0, 0) AND_177 (wire_525, {wire_526, wire_527});
or_n #(2, 0, 0) OR_83 (wire_528, {wire_395, wire_529});
notg #(0, 0) NOT_87 (wire_530, wire_383_11);
and_n #(2, 0, 0) AND_178 (wire_529, {wire_530, wire_531});
or_n #(2, 0, 0) OR_84 (wire_532, {wire_398, wire_533});
notg #(0, 0) NOT_88 (wire_534, wire_383_12);
and_n #(2, 0, 0) AND_179 (wire_533, {wire_534, wire_535});
or_n #(2, 0, 0) OR_85 (wire_536, {wire_401, wire_537});
notg #(0, 0) NOT_89 (wire_538, wire_383_13);
and_n #(2, 0, 0) AND_180 (wire_537, {wire_538, wire_539});
or_n #(2, 0, 0) OR_86 (wire_540, {wire_404, wire_541});
notg #(0, 0) NOT_90 (wire_542, wire_383_14);
and_n #(2, 0, 0) AND_181 (wire_541, {wire_542, wire_543});
nor_n #(2, 0, 0) NOR_2 (wire_383, {wire_457, wire_164});
or_n #(3, 0, 0) OR_87 (wire_544, {wire_27, wire_115, wire_164});
and_n #(2, 0, 0) AND_182 (wire_431, {wire_75, wire_545});
and_n #(2, 0, 0) AND_183 (wire_432, {wire_77, wire_546});
and_n #(2, 0, 0) AND_184 (wire_433, {wire_79, wire_547});
and_n #(2, 0, 0) AND_185 (wire_434, {wire_81, wire_548});
and_n #(2, 0, 0) AND_186 (wire_435, {wire_83, wire_549});
and_n #(2, 0, 0) AND_187 (wire_436, {wire_85, wire_550});
and_n #(2, 0, 0) AND_188 (wire_437, {wire_87, wire_551});
and_n #(2, 0, 0) AND_189 (wire_438, {wire_89, wire_552});
or_n #(2, 0, 0) OR_88 (wire_553, {wire_115, wire_164});
notg #(0, 0) NOT_91 (wire_554, wire_381);
notg #(0, 0) NOT_92 (wire_555, wire_556_0);
notg #(0, 0) NOT_93 (wire_557, wire_556_1);
notg #(0, 0) NOT_94 (wire_558, wire_556_2);
notg #(0, 0) NOT_95 (wire_559, wire_556_3);
notg #(0, 0) NOT_96 (wire_560, wire_556_4);
notg #(0, 0) NOT_97 (wire_561, wire_556_5);
notg #(0, 0) NOT_98 (wire_562, wire_556_6);
notg #(0, 0) NOT_99 (wire_563, wire_556_7);
notg #(0, 0) NOT_100 (wire_564, wire_556_8);
notg #(0, 0) NOT_101 (wire_565, wire_556_9);
notg #(0, 0) NOT_102 (wire_566, wire_556_10);
notg #(0, 0) NOT_103 (wire_567, wire_556_11);
notg #(0, 0) NOT_104 (wire_568, wire_556_12);
notg #(0, 0) NOT_105 (wire_569, wire_556_13);
notg #(0, 0) NOT_106 (wire_570, wire_556_14);
notg #(0, 0) NOT_107 (wire_571, wire_556_15);
notg #(0, 0) NOT_108 (wire_545, wire_556_16);
notg #(0, 0) NOT_109 (wire_546, wire_556_17);
notg #(0, 0) NOT_110 (wire_547, wire_556_18);
notg #(0, 0) NOT_111 (wire_548, wire_556_19);
notg #(0, 0) NOT_112 (wire_549, wire_556_20);
notg #(0, 0) NOT_113 (wire_550, wire_556_21);
notg #(0, 0) NOT_114 (wire_551, wire_556_22);
notg #(0, 0) NOT_115 (wire_552, wire_556_23);
notg #(0, 0) NOT_116 (wire_572, wire_556_24);
notg #(0, 0) NOT_117 (wire_573, wire_556_25);
notg #(0, 0) NOT_118 (wire_574, wire_556_26);
notg #(0, 0) NOT_119 (wire_575, wire_556_27);
notg #(0, 0) NOT_120 (wire_576, wire_556_28);
notg #(0, 0) NOT_121 (wire_577, wire_556_29);
notg #(0, 0) NOT_122 (wire_578, wire_556_30);
notg #(0, 0) NOT_123 (wire_579, wire_556_31);
notg #(0, 0) NOT_124 (wire_580, wire_556_32);
notg #(0, 0) NOT_125 (wire_581, wire_556_33);
notg #(0, 0) NOT_126 (wire_582, wire_556_34);
notg #(0, 0) NOT_127 (wire_583, wire_556_35);
notg #(0, 0) NOT_128 (wire_584, wire_556_36);
notg #(0, 0) NOT_129 (wire_585, wire_556_37);
notg #(0, 0) NOT_130 (wire_586, wire_556_38);
notg #(0, 0) NOT_131 (wire_587, wire_556_39);
notg #(0, 0) NOT_132 (wire_588, wire_556_40);
notg #(0, 0) NOT_133 (wire_589, wire_556_41);
notg #(0, 0) NOT_134 (wire_590, wire_556_42);
notg #(0, 0) NOT_135 (wire_591, wire_556_43);
notg #(0, 0) NOT_136 (wire_592, wire_556_44);
notg #(0, 0) NOT_137 (wire_593, wire_556_45);
notg #(0, 0) NOT_138 (wire_594, wire_556_46);
notg #(0, 0) NOT_139 (wire_595, wire_556_47);
notg #(0, 0) NOT_140 (wire_596, wire_556_48);
notg #(0, 0) NOT_141 (wire_597, wire_556_49);
notg #(0, 0) NOT_142 (wire_598, wire_556_50);
or_n #(2, 0, 0) OR_89 (wire_407, {wire_556_51, wire_381});
and_n #(2, 0, 0) AND_190 (wire_455, {wire_595, wire_457});
and_n #(2, 0, 0) AND_191 (wire_456, {wire_596, wire_27});
and_n #(2, 0, 0) AND_192 (wire_458, {wire_597, wire_115});
and_n #(2, 0, 0) AND_193 (wire_459, {wire_598, wire_164});
and_n #(2, 0, 0) AND_194 (wire_416, {wire_275, wire_579});
and_n #(2, 0, 0) AND_195 (wire_408, {wire_587, wire_324_1});
and_n #(2, 0, 0) AND_196 (wire_417, {wire_277, wire_580});
and_n #(2, 0, 0) AND_197 (wire_409, {wire_588, wire_326_1});
and_n #(2, 0, 0) AND_198 (wire_418, {wire_279, wire_581});
and_n #(2, 0, 0) AND_199 (wire_410, {wire_589, wire_328_1});
and_n #(2, 0, 0) AND_200 (wire_419, {wire_281, wire_582});
and_n #(2, 0, 0) AND_201 (wire_411, {wire_590, wire_330_1});
and_n #(2, 0, 0) AND_202 (wire_420, {wire_283, wire_583});
and_n #(2, 0, 0) AND_203 (wire_412, {wire_591, wire_332_1});
and_n #(2, 0, 0) AND_204 (wire_421, {wire_285, wire_584});
and_n #(2, 0, 0) AND_205 (wire_413, {wire_592, wire_334_1});
and_n #(2, 0, 0) AND_206 (wire_422, {wire_287, wire_585});
and_n #(2, 0, 0) AND_207 (wire_414, {wire_593, wire_336_1});
and_n #(2, 0, 0) AND_208 (wire_423, {wire_289, wire_586});
and_n #(2, 0, 0) AND_209 (wire_415, {wire_594, wire_338_1});
and_n #(2, 0, 0) AND_210 (wire_424, {wire_226, wire_572});
and_n #(2, 0, 0) AND_211 (wire_425, {wire_228, wire_573});
and_n #(2, 0, 0) AND_212 (wire_426, {wire_230, wire_574});
and_n #(2, 0, 0) AND_213 (wire_427, {wire_232, wire_575});
and_n #(2, 0, 0) AND_214 (wire_428, {wire_234, wire_576});
and_n #(2, 0, 0) AND_215 (wire_429, {wire_236, wire_577});
and_n #(2, 0, 0) AND_216 (wire_430, {wire_238, wire_578});
and_n #(2, 0, 0) AND_217 (wire_439, {wire_202, wire_564});
and_n #(2, 0, 0) AND_218 (wire_440, {wire_205, wire_565});
and_n #(2, 0, 0) AND_219 (wire_441, {wire_208, wire_566});
and_n #(2, 0, 0) AND_220 (wire_442, {wire_211, wire_567});
and_n #(2, 0, 0) AND_221 (wire_443, {wire_214, wire_568});
and_n #(2, 0, 0) AND_222 (wire_444, {wire_217, wire_569});
and_n #(2, 0, 0) AND_223 (wire_445, {wire_220, wire_570});
and_n #(2, 0, 0) AND_224 (wire_446, {wire_223, wire_571});
and_n #(2, 0, 0) AND_225 (wire_447, {wire_300, wire_555});
and_n #(2, 0, 0) AND_226 (wire_448, {wire_303, wire_557});
and_n #(2, 0, 0) AND_227 (wire_449, {wire_306, wire_558});
and_n #(2, 0, 0) AND_228 (wire_450, {wire_309, wire_559});
and_n #(2, 0, 0) AND_229 (wire_451, {wire_312, wire_560});
and_n #(2, 0, 0) AND_230 (wire_452, {wire_315, wire_561});
and_n #(2, 0, 0) AND_231 (wire_453, {wire_318, wire_562});
and_n #(2, 0, 0) AND_232 (wire_454, {wire_321, wire_563});
bufg #(0, 0) BUF_2 (wire_599, 1'b0);
notg #(0, 0) NOT_143 (wire_609, wire_556_52);
notg #(0, 0) NOT_144 (wire_610, wire_556_53);
notg #(0, 0) NOT_145 (wire_611, wire_556_54);
notg #(0, 0) NOT_146 (wire_612, wire_556_55);
notg #(0, 0) NOT_147 (wire_613, wire_556_56);
notg #(0, 0) NOT_148 (wire_614, wire_556_57);
notg #(0, 0) NOT_149 (wire_615, wire_556_58);
notg #(0, 0) NOT_150 (wire_616, wire_556_59);
and_n #(2, 0, 0) AND_233 (wire_601, {wire_382, wire_609});
and_n #(2, 0, 0) AND_234 (wire_602, {wire_516, wire_610});
and_n #(2, 0, 0) AND_235 (wire_603, {wire_520, wire_611});
and_n #(2, 0, 0) AND_236 (wire_604, {wire_524, wire_612});
and_n #(2, 0, 0) AND_237 (wire_605, {wire_528, wire_613});
and_n #(2, 0, 0) AND_238 (wire_606, {wire_532, wire_614});
and_n #(2, 0, 0) AND_239 (wire_607, {wire_536, wire_615});
and_n #(2, 0, 0) AND_240 (wire_608, {wire_540, wire_616});
bufg #(0, 0) BUF_3 (wire_600, 1'b1);
bufg #(0, 0) BUF_4 (wire_617, 1'b0);
or_n #(2, 0, 0) OR_90 (wire_618, {wire_554, wire_556_60});
notg #(0, 0) NOT_151 (wire_627, wire_556_61);
notg #(0, 0) NOT_152 (wire_628, wire_556_62);
notg #(0, 0) NOT_153 (wire_629, wire_556_63);
notg #(0, 0) NOT_154 (wire_630, wire_556_64);
notg #(0, 0) NOT_155 (wire_631, wire_556_65);
notg #(0, 0) NOT_156 (wire_632, wire_556_66);
notg #(0, 0) NOT_157 (wire_633, wire_556_67);
notg #(0, 0) NOT_158 (wire_634, wire_556_68);
and_n #(2, 0, 0) AND_241 (wire_619, {wire_491, wire_627});
and_n #(2, 0, 0) AND_242 (wire_620, {wire_495, wire_628});
and_n #(2, 0, 0) AND_243 (wire_621, {wire_498, wire_629});
and_n #(2, 0, 0) AND_244 (wire_622, {wire_501, wire_630});
and_n #(2, 0, 0) AND_245 (wire_623, {wire_504, wire_631});
and_n #(2, 0, 0) AND_246 (wire_624, {wire_507, wire_632});
and_n #(2, 0, 0) AND_247 (wire_625, {wire_510, wire_633});
and_n #(2, 0, 0) AND_248 (wire_626, {wire_513, wire_634});
bufg #(0, 0) BUF_5 (wire_635, 1'b0);
or_n #(2, 0, 0) OR_91 (wire_636, {wire_553, wire_556_69});
notg #(0, 0) NOT_159 (wire_645, wire_556_70);
notg #(0, 0) NOT_160 (wire_646, wire_556_71);
notg #(0, 0) NOT_161 (wire_647, wire_556_72);
notg #(0, 0) NOT_162 (wire_648, wire_556_73);
notg #(0, 0) NOT_163 (wire_649, wire_556_74);
notg #(0, 0) NOT_164 (wire_650, wire_556_75);
notg #(0, 0) NOT_165 (wire_651, wire_556_76);
notg #(0, 0) NOT_166 (wire_652, wire_556_77);
and_n #(2, 0, 0) AND_249 (wire_637, {wire_653, wire_645});
and_n #(2, 0, 0) AND_250 (wire_638, {wire_654, wire_646});
and_n #(2, 0, 0) AND_251 (wire_639, {wire_655, wire_647});
and_n #(2, 0, 0) AND_252 (wire_640, {wire_656, wire_648});
and_n #(2, 0, 0) AND_253 (wire_641, {wire_657, wire_649});
and_n #(2, 0, 0) AND_254 (wire_642, {wire_658, wire_650});
and_n #(2, 0, 0) AND_255 (wire_643, {wire_659, wire_651});
and_n #(2, 0, 0) AND_256 (wire_644, {wire_660, wire_652});
bufg #(0, 0) BUF_6 (wire_661, 1'b0);
or_n #(2, 0, 0) OR_92 (wire_662, {wire_544, wire_556_78});
notg #(0, 0) NOT_167 (wire_671, wire_556_79);
notg #(0, 0) NOT_168 (wire_672, wire_556_80);
notg #(0, 0) NOT_169 (wire_673, wire_556_81);
notg #(0, 0) NOT_170 (wire_674, wire_556_82);
notg #(0, 0) NOT_171 (wire_675, wire_556_83);
notg #(0, 0) NOT_172 (wire_676, wire_556_84);
notg #(0, 0) NOT_173 (wire_677, wire_556_85);
notg #(0, 0) NOT_174 (wire_678, wire_556_86);
and_n #(2, 0, 0) AND_257 (wire_663, {wire_460, wire_671});
and_n #(2, 0, 0) AND_258 (wire_664, {wire_463, wire_672});
and_n #(2, 0, 0) AND_259 (wire_665, {wire_467, wire_673});
and_n #(2, 0, 0) AND_260 (wire_666, {wire_471, wire_674});
and_n #(2, 0, 0) AND_261 (wire_667, {wire_475, wire_675});
and_n #(2, 0, 0) AND_262 (wire_668, {wire_479, wire_676});
and_n #(2, 0, 0) AND_263 (wire_669, {wire_483, wire_677});
and_n #(2, 0, 0) AND_264 (wire_670, {wire_487, wire_678});
xor_n #(2, 0, 0) XOR_1 (wire_523, {wire_679_0, wire_680_0});
xor_n #(2, 0, 0) XOR_2 (wire_681, {wire_682, wire_683});
xor_n #(2, 0, 0) XOR_3 (wire_682, {wire_684, wire_685});
xor_n #(2, 0, 0) XOR_4 (wire_686, {wire_687, wire_688_0});
xor_n #(2, 0, 0) XOR_5 (wire_687, {wire_689_0, wire_690_0});
xor_n #(2, 0, 0) XOR_6 (wire_691, {wire_692, wire_693_0});
xor_n #(2, 0, 0) XOR_7 (wire_692, {wire_694_0, wire_695_0});
xor_n #(2, 0, 0) XOR_8 (wire_696, {wire_697, wire_698_0});
xor_n #(2, 0, 0) XOR_9 (wire_697, {wire_699_0, wire_700_0});
xor_n #(2, 0, 0) XOR_10 (wire_701, {wire_702, wire_703_0});
xor_n #(2, 0, 0) XOR_11 (wire_702, {wire_704_0, wire_705_0});
bufg #(0, 0) BUF_7 (wire_680, wire_706);
and_n #(2, 0, 0) AND_265 (wire_703, {wire_680_1, wire_679_1});
bufg #(0, 0) BUF_8 (wire_704, wire_707);
and_n #(2, 0, 0) AND_266 (wire_708, {wire_704_1, wire_703_1});
or_n #(2, 0, 0) OR_93 (wire_709, {wire_704_2, wire_703_2});
bufg #(0, 0) BUF_9 (wire_699, wire_710);
and_n #(2, 0, 0) AND_267 (wire_711, {wire_699_1, wire_698_1});
or_n #(2, 0, 0) OR_94 (wire_712, {wire_699_2, wire_698_2});
bufg #(0, 0) BUF_10 (wire_694, wire_713);
and_n #(2, 0, 0) AND_268 (wire_714, {wire_694_1, wire_693_1});
or_n #(2, 0, 0) OR_95 (wire_715, {wire_694_2, wire_693_2});
bufg #(0, 0) BUF_11 (wire_689, wire_716);
and_n #(2, 0, 0) AND_269 (wire_717, {wire_689_1, wire_688_1});
or_n #(2, 0, 0) OR_96 (wire_718, {wire_689_2, wire_688_2});
bufg #(0, 0) BUF_12 (wire_684, wire_719);
bufg #(0, 0) BUF_13 (wire_527, wire_701);
bufg #(0, 0) BUF_14 (wire_720, wire_696);
bufg #(0, 0) BUF_15 (wire_721, wire_691);
bufg #(0, 0) BUF_16 (wire_722, wire_686);
bufg #(0, 0) BUF_17 (wire_723, wire_681);
bufg #(0, 0) BUF_18 (wire_531, wire_724);
bufg #(0, 0) BUF_19 (wire_724, wire_720);
bufg #(0, 0) BUF_20 (wire_725, wire_726);
bufg #(0, 0) BUF_21 (wire_726, wire_721);
bufg #(0, 0) BUF_22 (wire_727, wire_728);
bufg #(0, 0) BUF_23 (wire_728, wire_722);
bufg #(0, 0) BUF_24 (wire_729, wire_730);
bufg #(0, 0) BUF_25 (wire_730, wire_723);
bufg #(0, 0) BUF_26 (wire_535, wire_731);
bufg #(0, 0) BUF_27 (wire_731, wire_725);
bufg #(0, 0) BUF_28 (wire_732, wire_733);
bufg #(0, 0) BUF_29 (wire_733, wire_727);
bufg #(0, 0) BUF_30 (wire_734, wire_735);
bufg #(0, 0) BUF_31 (wire_735, wire_729);
bufg #(0, 0) BUF_32 (wire_539, wire_736);
bufg #(0, 0) BUF_33 (wire_736, wire_732);
bufg #(0, 0) BUF_34 (wire_737, wire_738);
bufg #(0, 0) BUF_35 (wire_738, wire_734);
bufg #(0, 0) BUF_36 (wire_543, wire_739);
bufg #(0, 0) BUF_37 (wire_739, wire_737);
bufg #(0, 0) BUF_38 (wire_706, wire_740);
bufg #(0, 0) BUF_39 (wire_707, wire_741);
bufg #(0, 0) BUF_40 (wire_710, wire_742);
bufg #(0, 0) BUF_41 (wire_713, wire_743);
bufg #(0, 0) BUF_42 (wire_716, wire_744);
bufg #(0, 0) BUF_43 (wire_719, wire_745);
and_n #(2, 0, 0) AND_270 (wire_745, {wire_199, wire_163_0});
and_n #(2, 0, 0) AND_271 (wire_744, {wire_198_0, wire_163_1});
and_n #(2, 0, 0) AND_272 (wire_743, {wire_197_0, wire_163_2});
and_n #(2, 0, 0) AND_273 (wire_742, {wire_196_0, wire_163_3});
and_n #(2, 0, 0) AND_274 (wire_741, {wire_195_0, wire_163_4});
and_n #(2, 0, 0) AND_275 (wire_740, {wire_194_0, wire_163_5});
bufg #(0, 0) BUF_44 (wire_519, wire_746);
and_n #(2, 0, 0) AND_276 (wire_746, {wire_193_0, wire_163_6});
and_n #(2, 0, 0) AND_277 (wire_685, {wire_198_1, wire_164});
and_n #(2, 0, 0) AND_278 (wire_690, {wire_197_1, wire_164});
and_n #(2, 0, 0) AND_279 (wire_747, {wire_690_1, wire_718});
and_n #(2, 0, 0) AND_280 (wire_695, {wire_196_1, wire_164});
and_n #(2, 0, 0) AND_281 (wire_748, {wire_695_1, wire_715});
and_n #(2, 0, 0) AND_282 (wire_700, {wire_195_1, wire_164});
and_n #(2, 0, 0) AND_283 (wire_749, {wire_700_1, wire_712});
and_n #(2, 0, 0) AND_284 (wire_705, {wire_194_1, wire_164});
and_n #(2, 0, 0) AND_285 (wire_750, {wire_705_1, wire_709});
and_n #(2, 0, 0) AND_286 (wire_679, {wire_193_1, wire_164});
or_n #(2, 0, 0) OR_97 (wire_698, {wire_708, wire_750});
or_n #(2, 0, 0) OR_98 (wire_693, {wire_711, wire_749});
or_n #(2, 0, 0) OR_99 (wire_688, {wire_714, wire_748});
or_n #(2, 0, 0) OR_100 (wire_683, {wire_717, wire_747});
xor_n #(2, 0, 0) XOR_12 (wire_497, {wire_751_0, wire_752_0});
xor_n #(2, 0, 0) XOR_13 (wire_500, {wire_753_0, wire_754_0});
xor_n #(2, 0, 0) XOR_14 (wire_755, {wire_756, wire_757});
xor_n #(2, 0, 0) XOR_15 (wire_756, {wire_758, wire_759});
xor_n #(2, 0, 0) XOR_16 (wire_760, {wire_761, wire_762_0});
xor_n #(2, 0, 0) XOR_17 (wire_761, {wire_763_0, wire_764_0});
xor_n #(2, 0, 0) XOR_18 (wire_765, {wire_766, wire_767_0});
xor_n #(2, 0, 0) XOR_19 (wire_766, {wire_768_0, wire_769_0});
xor_n #(2, 0, 0) XOR_20 (wire_770, {wire_771, wire_772_0});
xor_n #(2, 0, 0) XOR_21 (wire_771, {wire_773_0, wire_774_0});
xor_n #(2, 0, 0) XOR_22 (wire_775, {wire_776, wire_777_0});
xor_n #(2, 0, 0) XOR_23 (wire_776, {wire_778_0, wire_779_0});
xor_n #(2, 0, 0) XOR_24 (wire_758, {wire_780, wire_781});
xor_n #(2, 0, 0) XOR_25 (wire_780, {wire_782, wire_783});
xor_n #(2, 0, 0) XOR_26 (wire_763, {wire_784, wire_785_0});
xor_n #(2, 0, 0) XOR_27 (wire_784, {wire_786_0, wire_787_0});
xor_n #(2, 0, 0) XOR_28 (wire_768, {wire_788, wire_789_0});
xor_n #(2, 0, 0) XOR_29 (wire_788, {wire_790_0, wire_791_0});
xor_n #(2, 0, 0) XOR_30 (wire_773, {wire_792, wire_793_0});
xor_n #(2, 0, 0) XOR_31 (wire_792, {wire_794_0, wire_795_0});
xor_n #(2, 0, 0) XOR_32 (wire_778, {wire_796, wire_797_0});
xor_n #(2, 0, 0) XOR_33 (wire_796, {wire_798_0, wire_799_0});
xor_n #(2, 0, 0) XOR_34 (wire_754, {wire_800, wire_801_0});
xor_n #(2, 0, 0) XOR_35 (wire_800, {wire_802_0, wire_803_0});
and_n #(2, 0, 0) AND_287 (wire_777, {wire_754_1, wire_753_1});
and_n #(2, 0, 0) AND_288 (wire_804, {wire_778_1, wire_777_1});
or_n #(2, 0, 0) OR_101 (wire_805, {wire_778_2, wire_777_2});
and_n #(2, 0, 0) AND_289 (wire_806, {wire_773_1, wire_772_1});
or_n #(2, 0, 0) OR_102 (wire_807, {wire_773_2, wire_772_2});
and_n #(2, 0, 0) AND_290 (wire_808, {wire_768_1, wire_767_1});
or_n #(2, 0, 0) OR_103 (wire_809, {wire_768_2, wire_767_2});
and_n #(2, 0, 0) AND_291 (wire_810, {wire_763_1, wire_762_1});
or_n #(2, 0, 0) OR_104 (wire_811, {wire_763_2, wire_762_2});
bufg #(0, 0) BUF_45 (wire_503, wire_775);
bufg #(0, 0) BUF_46 (wire_812, wire_770);
bufg #(0, 0) BUF_47 (wire_813, wire_765);
bufg #(0, 0) BUF_48 (wire_814, wire_760);
bufg #(0, 0) BUF_49 (wire_815, wire_755);
bufg #(0, 0) BUF_50 (wire_506, wire_816);
bufg #(0, 0) BUF_51 (wire_816, wire_812);
bufg #(0, 0) BUF_52 (wire_817, wire_818);
bufg #(0, 0) BUF_53 (wire_818, wire_813);
bufg #(0, 0) BUF_54 (wire_819, wire_820);
bufg #(0, 0) BUF_55 (wire_820, wire_814);
bufg #(0, 0) BUF_56 (wire_821, wire_822);
bufg #(0, 0) BUF_57 (wire_822, wire_815);
bufg #(0, 0) BUF_58 (wire_509, wire_823);
bufg #(0, 0) BUF_59 (wire_823, wire_817);
bufg #(0, 0) BUF_60 (wire_824, wire_825);
bufg #(0, 0) BUF_61 (wire_825, wire_819);
bufg #(0, 0) BUF_62 (wire_826, wire_827);
bufg #(0, 0) BUF_63 (wire_827, wire_821);
bufg #(0, 0) BUF_64 (wire_512, wire_828);
bufg #(0, 0) BUF_65 (wire_828, wire_824);
bufg #(0, 0) BUF_66 (wire_829, wire_830);
bufg #(0, 0) BUF_67 (wire_830, wire_826);
bufg #(0, 0) BUF_68 (wire_515, wire_831);
bufg #(0, 0) BUF_69 (wire_831, wire_829);
and_n #(2, 0, 0) AND_292 (wire_782, {wire_248, wire_164});
and_n #(2, 0, 0) AND_293 (wire_832, {wire_786_1, wire_785_1});
and_n #(2, 0, 0) AND_294 (wire_833, {wire_786_2, wire_787_1});
and_n #(2, 0, 0) AND_295 (wire_786, {wire_247_0, wire_164});
and_n #(2, 0, 0) AND_296 (wire_790, {wire_246_0, wire_164});
and_n #(2, 0, 0) AND_297 (wire_834, {wire_790_1, wire_835});
and_n #(2, 0, 0) AND_298 (wire_794, {wire_245_0, wire_164});
and_n #(2, 0, 0) AND_299 (wire_836, {wire_794_1, wire_837});
and_n #(2, 0, 0) AND_300 (wire_798, {wire_244_0, wire_164});
and_n #(2, 0, 0) AND_301 (wire_838, {wire_798_1, wire_839});
and_n #(2, 0, 0) AND_302 (wire_802, {wire_243_0, wire_164});
and_n #(2, 0, 0) AND_303 (wire_840, {wire_802_1, wire_841});
and_n #(2, 0, 0) AND_304 (wire_801, {wire_752_1, wire_751_1});
and_n #(2, 0, 0) AND_305 (wire_752, {wire_242_0, wire_164});
and_n #(2, 0, 0) AND_306 (wire_783, {wire_247_1, wire_164});
and_n #(2, 0, 0) AND_307 (wire_842, {wire_787_2, wire_785_2});
and_n #(2, 0, 0) AND_308 (wire_787, {wire_246_1, wire_164});
and_n #(2, 0, 0) AND_309 (wire_791, {wire_245_1, wire_164});
and_n #(2, 0, 0) AND_310 (wire_843, {wire_791_1, wire_789_1});
or_n #(2, 0, 0) OR_105 (wire_835, {wire_791_2, wire_789_2});
and_n #(2, 0, 0) AND_311 (wire_795, {wire_244_1, wire_164});
and_n #(2, 0, 0) AND_312 (wire_844, {wire_795_1, wire_793_1});
or_n #(2, 0, 0) OR_106 (wire_837, {wire_795_2, wire_793_2});
and_n #(2, 0, 0) AND_313 (wire_799, {wire_243_1, wire_164});
and_n #(2, 0, 0) AND_314 (wire_845, {wire_799_1, wire_797_1});
or_n #(2, 0, 0) OR_107 (wire_839, {wire_799_2, wire_797_2});
and_n #(2, 0, 0) AND_315 (wire_803, {wire_242_1, wire_164});
and_n #(2, 0, 0) AND_316 (wire_846, {wire_803_1, wire_801_1});
or_n #(2, 0, 0) OR_108 (wire_841, {wire_803_2, wire_801_2});
and_n #(2, 0, 0) AND_317 (wire_751, {wire_241_0, wire_164});
and_n #(2, 0, 0) AND_318 (wire_759, {wire_246_2, wire_200_0});
and_n #(2, 0, 0) AND_319 (wire_764, {wire_245_2, wire_200_1});
and_n #(2, 0, 0) AND_320 (wire_847, {wire_764_1, wire_811});
and_n #(2, 0, 0) AND_321 (wire_769, {wire_244_2, wire_200_2});
and_n #(2, 0, 0) AND_322 (wire_848, {wire_769_1, wire_809});
and_n #(2, 0, 0) AND_323 (wire_774, {wire_243_2, wire_200_3});
and_n #(2, 0, 0) AND_324 (wire_849, {wire_774_1, wire_807});
and_n #(2, 0, 0) AND_325 (wire_779, {wire_242_2, wire_200_4});
and_n #(2, 0, 0) AND_326 (wire_850, {wire_779_1, wire_805});
and_n #(2, 0, 0) AND_327 (wire_753, {wire_241_1, wire_200_5});
or_n #(2, 0, 0) OR_109 (wire_797, {wire_846, wire_840});
or_n #(2, 0, 0) OR_110 (wire_793, {wire_845, wire_838});
or_n #(2, 0, 0) OR_111 (wire_789, {wire_844, wire_836});
or_n #(2, 0, 0) OR_112 (wire_785, {wire_843, wire_834});
or_n #(3, 0, 0) OR_113 (wire_781, {wire_833, wire_832, wire_842});
or_n #(2, 0, 0) OR_114 (wire_772, {wire_804, wire_850});
or_n #(2, 0, 0) OR_115 (wire_767, {wire_806, wire_849});
or_n #(2, 0, 0) OR_116 (wire_762, {wire_808, wire_848});
or_n #(2, 0, 0) OR_117 (wire_757, {wire_810, wire_847});
and_n #(2, 0, 0) AND_328 (wire_494, {wire_241_2, wire_164});
xor_n #(2, 0, 0) XOR_36 (wire_654, {wire_290_0, wire_851_0});
xor_n #(2, 0, 0) XOR_37 (wire_852, {wire_853, wire_854});
xor_n #(2, 0, 0) XOR_38 (wire_853, {wire_855, wire_296_0});
xor_n #(2, 0, 0) XOR_39 (wire_856, {wire_857, wire_858_0});
xor_n #(2, 0, 0) XOR_40 (wire_857, {wire_859_0, wire_295_0});
xor_n #(2, 0, 0) XOR_41 (wire_860, {wire_861, wire_862_0});
xor_n #(2, 0, 0) XOR_42 (wire_861, {wire_863_0, wire_294_0});
xor_n #(2, 0, 0) XOR_43 (wire_864, {wire_865, wire_866_0});
xor_n #(2, 0, 0) XOR_44 (wire_865, {wire_867_0, wire_293_0});
xor_n #(2, 0, 0) XOR_45 (wire_868, {wire_869, wire_870_0});
xor_n #(2, 0, 0) XOR_46 (wire_869, {wire_871_0, wire_292_0});
xor_n #(2, 0, 0) XOR_47 (wire_872, {wire_873, wire_874_0});
xor_n #(2, 0, 0) XOR_48 (wire_873, {wire_875_0, wire_291_0});
bufg #(0, 0) BUF_70 (wire_655, wire_872);
bufg #(0, 0) BUF_71 (wire_876, wire_868);
bufg #(0, 0) BUF_72 (wire_877, wire_864);
bufg #(0, 0) BUF_73 (wire_878, wire_860);
bufg #(0, 0) BUF_74 (wire_879, wire_856);
bufg #(0, 0) BUF_75 (wire_880, wire_852);
bufg #(0, 0) BUF_76 (wire_656, wire_881);
bufg #(0, 0) BUF_77 (wire_881, wire_876);
bufg #(0, 0) BUF_78 (wire_882, wire_883);
bufg #(0, 0) BUF_79 (wire_883, wire_877);
bufg #(0, 0) BUF_80 (wire_884, wire_885);
bufg #(0, 0) BUF_81 (wire_885, wire_878);
bufg #(0, 0) BUF_82 (wire_886, wire_887);
bufg #(0, 0) BUF_83 (wire_887, wire_879);
bufg #(0, 0) BUF_84 (wire_888, wire_889);
bufg #(0, 0) BUF_85 (wire_889, wire_880);
bufg #(0, 0) BUF_86 (wire_657, wire_890);
bufg #(0, 0) BUF_87 (wire_890, wire_882);
bufg #(0, 0) BUF_88 (wire_891, wire_892);
bufg #(0, 0) BUF_89 (wire_892, wire_884);
bufg #(0, 0) BUF_90 (wire_893, wire_894);
bufg #(0, 0) BUF_91 (wire_894, wire_886);
bufg #(0, 0) BUF_92 (wire_895, wire_896);
bufg #(0, 0) BUF_93 (wire_896, wire_888);
bufg #(0, 0) BUF_94 (wire_658, wire_897);
bufg #(0, 0) BUF_95 (wire_897, wire_891);
bufg #(0, 0) BUF_96 (wire_898, wire_899);
bufg #(0, 0) BUF_97 (wire_899, wire_893);
bufg #(0, 0) BUF_98 (wire_900, wire_901);
bufg #(0, 0) BUF_99 (wire_901, wire_895);
bufg #(0, 0) BUF_100 (wire_659, wire_902);
bufg #(0, 0) BUF_101 (wire_902, wire_898);
bufg #(0, 0) BUF_102 (wire_903, wire_904);
bufg #(0, 0) BUF_103 (wire_904, wire_900);
bufg #(0, 0) BUF_104 (wire_660, wire_905);
bufg #(0, 0) BUF_105 (wire_905, wire_903);
and_n #(2, 0, 0) AND_329 (wire_855, {wire_297, wire_249_0});
and_n #(2, 0, 0) AND_330 (wire_906, {wire_859_1, wire_858_1});
and_n #(2, 0, 0) AND_331 (wire_907, {wire_859_2, wire_295_1});
and_n #(2, 0, 0) AND_332 (wire_859, {wire_296_1, wire_249_1});
and_n #(2, 0, 0) AND_333 (wire_863, {wire_295_2, wire_249_2});
and_n #(2, 0, 0) AND_334 (wire_908, {wire_863_1, wire_909});
and_n #(2, 0, 0) AND_335 (wire_867, {wire_294_1, wire_249_3});
and_n #(2, 0, 0) AND_336 (wire_910, {wire_867_1, wire_911});
and_n #(2, 0, 0) AND_337 (wire_871, {wire_293_1, wire_249_4});
and_n #(2, 0, 0) AND_338 (wire_912, {wire_871_1, wire_913});
and_n #(2, 0, 0) AND_339 (wire_875, {wire_292_1, wire_249_5});
and_n #(2, 0, 0) AND_340 (wire_914, {wire_875_1, wire_915});
and_n #(2, 0, 0) AND_341 (wire_874, {wire_851_1, wire_290_1});
and_n #(2, 0, 0) AND_342 (wire_851, {wire_291_1, wire_249_6});
and_n #(2, 0, 0) AND_343 (wire_916, {wire_874_1, wire_291_2});
or_n #(2, 0, 0) OR_118 (wire_915, {wire_874_2, wire_291_3});
or_n #(2, 0, 0) OR_119 (wire_870, {wire_916, wire_914});
and_n #(2, 0, 0) AND_344 (wire_917, {wire_870_1, wire_292_2});
or_n #(2, 0, 0) OR_120 (wire_913, {wire_870_2, wire_292_3});
or_n #(2, 0, 0) OR_121 (wire_866, {wire_917, wire_912});
and_n #(2, 0, 0) AND_345 (wire_918, {wire_866_1, wire_293_2});
or_n #(2, 0, 0) OR_122 (wire_911, {wire_866_2, wire_293_3});
or_n #(2, 0, 0) OR_123 (wire_862, {wire_918, wire_910});
and_n #(2, 0, 0) AND_346 (wire_919, {wire_862_1, wire_294_2});
or_n #(2, 0, 0) OR_124 (wire_909, {wire_862_2, wire_294_3});
and_n #(2, 0, 0) AND_347 (wire_920, {wire_858_2, wire_295_3});
or_n #(2, 0, 0) OR_125 (wire_858, {wire_919, wire_908});
or_n #(3, 0, 0) OR_126 (wire_854, {wire_907, wire_906, wire_920});
and_n #(2, 0, 0) AND_348 (wire_653, {wire_290_2, wire_249_7});
xor_n #(2, 0, 0) XOR_49 (wire_466, {wire_921_0, wire_340_0});
xor_n #(2, 0, 0) XOR_50 (wire_470, {wire_922_0, wire_923_0});
xor_n #(2, 0, 0) XOR_51 (wire_924, {wire_925, wire_926});
xor_n #(2, 0, 0) XOR_52 (wire_925, {wire_927, wire_928});
xor_n #(2, 0, 0) XOR_53 (wire_929, {wire_930, wire_931_0});
xor_n #(2, 0, 0) XOR_54 (wire_930, {wire_932_0, wire_933_0});
xor_n #(2, 0, 0) XOR_55 (wire_934, {wire_935, wire_936_0});
xor_n #(2, 0, 0) XOR_56 (wire_935, {wire_937_0, wire_938_0});
xor_n #(2, 0, 0) XOR_57 (wire_939, {wire_940, wire_941_0});
xor_n #(2, 0, 0) XOR_58 (wire_940, {wire_942_0, wire_943_0});
xor_n #(2, 0, 0) XOR_59 (wire_944, {wire_945, wire_946_0});
xor_n #(2, 0, 0) XOR_60 (wire_945, {wire_947_0, wire_948_0});
xor_n #(2, 0, 0) XOR_61 (wire_927, {wire_949, wire_950});
xor_n #(2, 0, 0) XOR_62 (wire_949, {wire_346, wire_951});
xor_n #(2, 0, 0) XOR_63 (wire_932, {wire_952, wire_953_0});
xor_n #(2, 0, 0) XOR_64 (wire_952, {wire_345_0, wire_954_0});
xor_n #(2, 0, 0) XOR_65 (wire_937, {wire_955, wire_956_0});
xor_n #(2, 0, 0) XOR_66 (wire_955, {wire_344_0, wire_957_0});
xor_n #(2, 0, 0) XOR_67 (wire_942, {wire_958, wire_959_0});
xor_n #(2, 0, 0) XOR_68 (wire_958, {wire_343_0, wire_960_0});
xor_n #(2, 0, 0) XOR_69 (wire_947, {wire_961, wire_962_0});
xor_n #(2, 0, 0) XOR_70 (wire_961, {wire_342_0, wire_963_0});
xor_n #(2, 0, 0) XOR_71 (wire_923, {wire_964, wire_965_0});
xor_n #(2, 0, 0) XOR_72 (wire_964, {wire_341_0, wire_966_0});
and_n #(2, 0, 0) AND_349 (wire_946, {wire_923_1, wire_922_1});
and_n #(2, 0, 0) AND_350 (wire_967, {wire_947_1, wire_946_1});
or_n #(2, 0, 0) OR_127 (wire_968, {wire_947_2, wire_946_2});
and_n #(2, 0, 0) AND_351 (wire_969, {wire_942_1, wire_941_1});
or_n #(2, 0, 0) OR_128 (wire_970, {wire_942_2, wire_941_2});
and_n #(2, 0, 0) AND_352 (wire_971, {wire_937_1, wire_936_1});
or_n #(2, 0, 0) OR_129 (wire_972, {wire_937_2, wire_936_2});
and_n #(2, 0, 0) AND_353 (wire_973, {wire_932_1, wire_931_1});
or_n #(2, 0, 0) OR_130 (wire_974, {wire_932_2, wire_931_2});
bufg #(0, 0) BUF_106 (wire_474, wire_944);
bufg #(0, 0) BUF_107 (wire_975, wire_939);
bufg #(0, 0) BUF_108 (wire_976, wire_934);
bufg #(0, 0) BUF_109 (wire_977, wire_929);
bufg #(0, 0) BUF_110 (wire_978, wire_924);
bufg #(0, 0) BUF_111 (wire_478, wire_979);
bufg #(0, 0) BUF_112 (wire_979, wire_975);
bufg #(0, 0) BUF_113 (wire_980, wire_981);
bufg #(0, 0) BUF_114 (wire_981, wire_976);
bufg #(0, 0) BUF_115 (wire_982, wire_983);
bufg #(0, 0) BUF_116 (wire_983, wire_977);
bufg #(0, 0) BUF_117 (wire_984, wire_985);
bufg #(0, 0) BUF_118 (wire_985, wire_978);
bufg #(0, 0) BUF_119 (wire_482, wire_986);
bufg #(0, 0) BUF_120 (wire_986, wire_980);
bufg #(0, 0) BUF_121 (wire_987, wire_988);
bufg #(0, 0) BUF_122 (wire_988, wire_982);
bufg #(0, 0) BUF_123 (wire_989, wire_990);
bufg #(0, 0) BUF_124 (wire_990, wire_984);
bufg #(0, 0) BUF_125 (wire_486, wire_991);
bufg #(0, 0) BUF_126 (wire_991, wire_987);
bufg #(0, 0) BUF_127 (wire_992, wire_993);
bufg #(0, 0) BUF_128 (wire_993, wire_989);
bufg #(0, 0) BUF_129 (wire_490, wire_994);
bufg #(0, 0) BUF_130 (wire_994, wire_992);
and_n #(2, 0, 0) AND_354 (wire_951, {wire_345_1, wire_164});
and_n #(2, 0, 0) AND_355 (wire_995, {wire_954_1, wire_953_1});
and_n #(2, 0, 0) AND_356 (wire_996, {wire_954_2, wire_345_2});
and_n #(2, 0, 0) AND_357 (wire_954, {wire_344_1, wire_164});
and_n #(2, 0, 0) AND_358 (wire_957, {wire_343_1, wire_164});
and_n #(2, 0, 0) AND_359 (wire_997, {wire_957_1, wire_956_1});
or_n #(2, 0, 0) OR_131 (wire_998, {wire_957_2, wire_956_2});
and_n #(2, 0, 0) AND_360 (wire_960, {wire_342_1, wire_164});
and_n #(2, 0, 0) AND_361 (wire_999, {wire_960_1, wire_959_1});
or_n #(2, 0, 0) OR_132 (wire_1000, {wire_960_2, wire_959_2});
and_n #(2, 0, 0) AND_362 (wire_963, {wire_341_1, wire_164});
and_n #(2, 0, 0) AND_363 (wire_1001, {wire_963_1, wire_962_1});
or_n #(2, 0, 0) OR_133 (wire_1002, {wire_963_2, wire_962_2});
and_n #(2, 0, 0) AND_364 (wire_966, {wire_340_1, wire_164});
and_n #(2, 0, 0) AND_365 (wire_1003, {wire_966_1, wire_965_1});
or_n #(2, 0, 0) OR_134 (wire_1004, {wire_966_2, wire_965_2});
and_n #(2, 0, 0) AND_366 (wire_965, {wire_921_1, wire_340_2});
and_n #(2, 0, 0) AND_367 (wire_921, {wire_164, wire_339_1});
and_n #(2, 0, 0) AND_368 (wire_928, {wire_344_2, wire_298_0});
and_n #(2, 0, 0) AND_369 (wire_933, {wire_343_2, wire_298_1});
and_n #(2, 0, 0) AND_370 (wire_1005, {wire_933_1, wire_974});
and_n #(2, 0, 0) AND_371 (wire_938, {wire_342_2, wire_298_2});
and_n #(2, 0, 0) AND_372 (wire_1006, {wire_938_1, wire_972});
and_n #(2, 0, 0) AND_373 (wire_943, {wire_341_2, wire_298_3});
and_n #(2, 0, 0) AND_374 (wire_1007, {wire_943_1, wire_970});
and_n #(2, 0, 0) AND_375 (wire_948, {wire_340_3, wire_298_4});
and_n #(2, 0, 0) AND_376 (wire_1008, {wire_948_1, wire_968});
and_n #(2, 0, 0) AND_377 (wire_922, {wire_298_5, wire_339_2});
or_n #(2, 0, 0) OR_135 (wire_962, {wire_1003, wire_1009});
and_n #(2, 0, 0) AND_378 (wire_1009, {wire_1004, wire_341_3});
or_n #(2, 0, 0) OR_136 (wire_959, {wire_1001, wire_1010});
and_n #(2, 0, 0) AND_379 (wire_1010, {wire_1002, wire_342_3});
or_n #(2, 0, 0) OR_137 (wire_956, {wire_999, wire_1011});
and_n #(2, 0, 0) AND_380 (wire_1011, {wire_1000, wire_343_3});
and_n #(2, 0, 0) AND_381 (wire_1012, {wire_953_2, wire_345_3});
or_n #(2, 0, 0) OR_138 (wire_953, {wire_997, wire_1013});
and_n #(2, 0, 0) AND_382 (wire_1013, {wire_998, wire_344_3});
or_n #(3, 0, 0) OR_139 (wire_950, {wire_996, wire_1012, wire_995});
or_n #(2, 0, 0) OR_140 (wire_941, {wire_967, wire_1008});
or_n #(2, 0, 0) OR_141 (wire_936, {wire_969, wire_1007});
or_n #(2, 0, 0) OR_142 (wire_931, {wire_971, wire_1006});
or_n #(2, 0, 0) OR_143 (wire_926, {wire_973, wire_1005});
xor_n #(2, 0, 0) XOR_73 (wire_380, {wire_42_0, wire_90_0});
xor_n #(2, 0, 0) XOR_74 (wire_403, {wire_1014, wire_1015});
xor_n #(2, 0, 0) XOR_75 (wire_1014, {wire_97, wire_49});
xor_n #(2, 0, 0) XOR_76 (wire_400, {wire_1016, wire_1017_0});
xor_n #(2, 0, 0) XOR_77 (wire_1016, {wire_96_0, wire_48_0});
xor_n #(2, 0, 0) XOR_78 (wire_397, {wire_1018, wire_1019_0});
xor_n #(2, 0, 0) XOR_79 (wire_1018, {wire_95_0, wire_47_0});
xor_n #(2, 0, 0) XOR_80 (wire_394, {wire_1020, wire_1021_0});
xor_n #(2, 0, 0) XOR_81 (wire_1020, {wire_94_0, wire_46_0});
xor_n #(2, 0, 0) XOR_82 (wire_391, {wire_1022, wire_1023_0});
xor_n #(2, 0, 0) XOR_83 (wire_1022, {wire_93_0, wire_45_0});
xor_n #(2, 0, 0) XOR_84 (wire_388, {wire_1024, wire_1025_0});
xor_n #(2, 0, 0) XOR_85 (wire_1024, {wire_92_0, wire_44_0});
xor_n #(2, 0, 0) XOR_86 (wire_385, {wire_1026, wire_1027_0});
xor_n #(2, 0, 0) XOR_87 (wire_1026, {wire_91_0, wire_43_0});
and_n #(2, 0, 0) AND_383 (wire_1027, {wire_90_1, wire_42_1});
and_n #(2, 0, 0) AND_384 (wire_1028, {wire_1027_1, wire_43_1});
or_n #(2, 0, 0) OR_144 (wire_1029, {wire_1027_2, wire_43_2});
or_n #(2, 0, 0) OR_145 (wire_1025, {wire_1028, wire_1030});
and_n #(2, 0, 0) AND_385 (wire_1031, {wire_1025_1, wire_44_1});
or_n #(2, 0, 0) OR_146 (wire_1032, {wire_1025_2, wire_44_2});
and_n #(2, 0, 0) AND_386 (wire_1030, {wire_1029, wire_91_1});
or_n #(2, 0, 0) OR_147 (wire_1023, {wire_1031, wire_1033});
and_n #(2, 0, 0) AND_387 (wire_1034, {wire_1023_1, wire_45_1});
or_n #(2, 0, 0) OR_148 (wire_1035, {wire_1023_2, wire_45_2});
and_n #(2, 0, 0) AND_388 (wire_1033, {wire_1032, wire_92_1});
or_n #(2, 0, 0) OR_149 (wire_1021, {wire_1034, wire_1036});
and_n #(2, 0, 0) AND_389 (wire_1037, {wire_1021_1, wire_46_1});
or_n #(2, 0, 0) OR_150 (wire_1038, {wire_1021_2, wire_46_2});
and_n #(2, 0, 0) AND_390 (wire_1036, {wire_1035, wire_93_1});
or_n #(2, 0, 0) OR_151 (wire_1019, {wire_1037, wire_1039});
and_n #(2, 0, 0) AND_391 (wire_1040, {wire_1019_1, wire_47_1});
or_n #(2, 0, 0) OR_152 (wire_1041, {wire_1019_2, wire_47_2});
and_n #(2, 0, 0) AND_392 (wire_1039, {wire_1038, wire_94_1});
and_n #(2, 0, 0) AND_393 (wire_1042, {wire_1017_1, wire_48_1});
and_n #(2, 0, 0) AND_394 (wire_1043, {wire_1017_2, wire_96_1});
or_n #(2, 0, 0) OR_153 (wire_1017, {wire_1040, wire_1044});
and_n #(2, 0, 0) AND_395 (wire_1044, {wire_1041, wire_95_1});
or_n #(3, 0, 0) OR_154 (wire_1015, {wire_1045, wire_1043, wire_1042});
and_n #(2, 0, 0) AND_396 (wire_1045, {wire_96_2, wire_48_2});
xor_n #(2, 0, 0) XOR_88 (wire_348, {wire_123_0, wire_155_0});
xor_n #(2, 0, 0) XOR_89 (wire_376, {wire_1046, wire_1047});
xor_n #(2, 0, 0) XOR_90 (wire_1046, {wire_162, wire_130});
xor_n #(2, 0, 0) XOR_91 (wire_372, {wire_1048, wire_1049_0});
xor_n #(2, 0, 0) XOR_92 (wire_1048, {wire_161_0, wire_129_0});
xor_n #(2, 0, 0) XOR_93 (wire_368, {wire_1050, wire_1051_0});
xor_n #(2, 0, 0) XOR_94 (wire_1050, {wire_160_0, wire_128_0});
xor_n #(2, 0, 0) XOR_95 (wire_364, {wire_1052, wire_1053_0});
xor_n #(2, 0, 0) XOR_96 (wire_1052, {wire_159_0, wire_127_0});
xor_n #(2, 0, 0) XOR_97 (wire_360, {wire_1054, wire_1055_0});
xor_n #(2, 0, 0) XOR_98 (wire_1054, {wire_158_0, wire_126_0});
xor_n #(2, 0, 0) XOR_99 (wire_356, {wire_1056, wire_1057_0});
xor_n #(2, 0, 0) XOR_100 (wire_1056, {wire_157_0, wire_125_0});
xor_n #(2, 0, 0) XOR_101 (wire_352, {wire_1058, wire_1059_0});
xor_n #(2, 0, 0) XOR_102 (wire_1058, {wire_156_0, wire_124_0});
and_n #(2, 0, 0) AND_397 (wire_1059, {wire_155_1, wire_123_1});
and_n #(2, 0, 0) AND_398 (wire_1060, {wire_1059_1, wire_124_1});
or_n #(2, 0, 0) OR_155 (wire_1061, {wire_1059_2, wire_124_2});
or_n #(2, 0, 0) OR_156 (wire_1057, {wire_1060, wire_1062});
and_n #(2, 0, 0) AND_399 (wire_1063, {wire_1057_1, wire_125_1});
or_n #(2, 0, 0) OR_157 (wire_1064, {wire_1057_2, wire_125_2});
and_n #(2, 0, 0) AND_400 (wire_1062, {wire_1061, wire_156_1});
or_n #(2, 0, 0) OR_158 (wire_1055, {wire_1063, wire_1065});
and_n #(2, 0, 0) AND_401 (wire_1066, {wire_1055_1, wire_126_1});
or_n #(2, 0, 0) OR_159 (wire_1067, {wire_1055_2, wire_126_2});
and_n #(2, 0, 0) AND_402 (wire_1065, {wire_1064, wire_157_1});
or_n #(2, 0, 0) OR_160 (wire_1053, {wire_1066, wire_1068});
and_n #(2, 0, 0) AND_403 (wire_1069, {wire_1053_1, wire_127_1});
or_n #(2, 0, 0) OR_161 (wire_1070, {wire_1053_2, wire_127_2});
and_n #(2, 0, 0) AND_404 (wire_1068, {wire_1067, wire_158_1});
or_n #(2, 0, 0) OR_162 (wire_1051, {wire_1069, wire_1071});
and_n #(2, 0, 0) AND_405 (wire_1072, {wire_1051_1, wire_128_1});
or_n #(2, 0, 0) OR_163 (wire_1073, {wire_1051_2, wire_128_2});
and_n #(2, 0, 0) AND_406 (wire_1071, {wire_1070, wire_159_1});
and_n #(2, 0, 0) AND_407 (wire_1074, {wire_1049_1, wire_129_1});
and_n #(2, 0, 0) AND_408 (wire_1075, {wire_1049_2, wire_161_1});
or_n #(2, 0, 0) OR_164 (wire_1049, {wire_1072, wire_1076});
and_n #(2, 0, 0) AND_409 (wire_1076, {wire_1073, wire_160_1});
or_n #(3, 0, 0) OR_165 (wire_1047, {wire_1077, wire_1075, wire_1074});
and_n #(2, 0, 0) AND_410 (wire_1077, {wire_161_2, wire_129_2});
bufg #(0, 0) BUF_131 (wire_406, clk_net_0);
bufg #(0, 0) BUF_132 (wire_556, reset_net_0);
bufg #(0, 0) BUF_133 (wire_324, x_7);
bufg #(0, 0) BUF_134 (wire_326, x_6);
bufg #(0, 0) BUF_135 (wire_328, x_5);
bufg #(0, 0) BUF_136 (wire_330, x_4);
bufg #(0, 0) BUF_137 (wire_332, x_3);
bufg #(0, 0) BUF_138 (wire_334, x_2);
bufg #(0, 0) BUF_139 (wire_336, x_1);
bufg #(0, 0) BUF_140 (wire_338, x_0);
bufg #(0, 0) BUF_141 (y_7, wire_379);
bufg #(0, 0) BUF_142 (y_6, wire_384);
bufg #(0, 0) BUF_143 (y_5, wire_387);
bufg #(0, 0) BUF_144 (y_4, wire_390);
bufg #(0, 0) BUF_145 (y_3, wire_393);
bufg #(0, 0) BUF_146 (y_2, wire_396);
bufg #(0, 0) BUF_147 (y_1, wire_399);
bufg #(0, 0) BUF_148 (y_0, wire_402);
dff DFF_1  (wire_275, wire_408, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_2  (wire_277, wire_409, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_3  (wire_279, wire_410, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_4  (wire_281, wire_411, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_5  (wire_283, wire_412, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_6  (wire_285, wire_413, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_7  (wire_287, wire_414, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_8  (wire_289, wire_415, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_9  (wire_226, wire_416, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_10  (wire_228, wire_417, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_11  (wire_230, wire_418, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_12  (wire_232, wire_419, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_13  (wire_234, wire_420, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_14  (wire_236, wire_421, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_15  (wire_238, wire_422, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_16  (wire_240, wire_423, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_17  (wire_180, wire_424, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_18  (wire_182, wire_425, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_19  (wire_184, wire_426, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_20  (wire_186, wire_427, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_21  (wire_188, wire_428, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_22  (wire_190, wire_429, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_23  (wire_192, wire_430, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_24  (wire_202, wire_431, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_25  (wire_205, wire_432, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_26  (wire_208, wire_433, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_27  (wire_211, wire_434, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_28  (wire_214, wire_435, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_29  (wire_217, wire_436, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_30  (wire_220, wire_437, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_31  (wire_223, wire_438, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_32  (wire_300, wire_439, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_33  (wire_303, wire_440, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_34  (wire_306, wire_441, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_35  (wire_309, wire_442, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_36  (wire_312, wire_443, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_37  (wire_315, wire_444, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_38  (wire_318, wire_445, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_39  (wire_321, wire_446, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_40  (wire_251, wire_447, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_41  (wire_254, wire_448, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_42  (wire_257, wire_449, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_43  (wire_260, wire_450, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_44  (wire_263, wire_451, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_45  (wire_266, wire_452, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_46  (wire_269, wire_453, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_47  (wire_272, wire_454, wire_406, wire_405, 1'b0, wire_407, NbarT, Si, 1'b0);
dff DFF_48  (wire_381, wire_455, wire_406, 1'b0, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_49  (wire_457, wire_456, wire_406, 1'b0, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_50  (wire_27, wire_458, wire_406, 1'b0, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_51  (wire_115, wire_459, wire_406, 1'b0, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_52  (wire_164, wire_407, wire_406, 1'b0, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_53  (wire_2, wire_601, wire_406, wire_599, 1'b0, wire_600, NbarT, Si, 1'b0);
dff DFF_54  (wire_5, wire_602, wire_406, wire_599, 1'b0, wire_600, NbarT, Si, 1'b0);
dff DFF_55  (wire_8, wire_603, wire_406, wire_599, 1'b0, wire_600, NbarT, Si, 1'b0);
dff DFF_56  (wire_11, wire_604, wire_406, wire_599, 1'b0, wire_600, NbarT, Si, 1'b0);
dff DFF_57  (wire_14, wire_605, wire_406, wire_599, 1'b0, wire_600, NbarT, Si, 1'b0);
dff DFF_58  (wire_17, wire_606, wire_406, wire_599, 1'b0, wire_600, NbarT, Si, 1'b0);
dff DFF_59  (wire_20, wire_607, wire_406, wire_599, 1'b0, wire_600, NbarT, Si, 1'b0);
dff DFF_60  (wire_23, wire_608, wire_406, wire_599, 1'b0, wire_600, NbarT, Si, 1'b0);
dff DFF_61  (wire_51, wire_619, wire_406, wire_617, 1'b0, wire_618, NbarT, Si, 1'b0);
dff DFF_62  (wire_54, wire_620, wire_406, wire_617, 1'b0, wire_618, NbarT, Si, 1'b0);
dff DFF_63  (wire_57, wire_621, wire_406, wire_617, 1'b0, wire_618, NbarT, Si, 1'b0);
dff DFF_64  (wire_60, wire_622, wire_406, wire_617, 1'b0, wire_618, NbarT, Si, 1'b0);
dff DFF_65  (wire_63, wire_623, wire_406, wire_617, 1'b0, wire_618, NbarT, Si, 1'b0);
dff DFF_66  (wire_66, wire_624, wire_406, wire_617, 1'b0, wire_618, NbarT, Si, 1'b0);
dff DFF_67  (wire_69, wire_625, wire_406, wire_617, 1'b0, wire_618, NbarT, Si, 1'b0);
dff DFF_68  (wire_72, wire_626, wire_406, wire_617, 1'b0, wire_618, NbarT, Si, 1'b0);
dff DFF_69  (wire_26, wire_637, wire_406, wire_635, 1'b0, wire_636, NbarT, Si, 1'b0);
dff DFF_70  (wire_29, wire_638, wire_406, wire_635, 1'b0, wire_636, NbarT, Si, 1'b0);
dff DFF_71  (wire_31, wire_639, wire_406, wire_635, 1'b0, wire_636, NbarT, Si, 1'b0);
dff DFF_72  (wire_33, wire_640, wire_406, wire_635, 1'b0, wire_636, NbarT, Si, 1'b0);
dff DFF_73  (wire_35, wire_641, wire_406, wire_635, 1'b0, wire_636, NbarT, Si, 1'b0);
dff DFF_74  (wire_37, wire_642, wire_406, wire_635, 1'b0, wire_636, NbarT, Si, 1'b0);
dff DFF_75  (wire_39, wire_643, wire_406, wire_635, 1'b0, wire_636, NbarT, Si, 1'b0);
dff DFF_76  (wire_41, wire_644, wire_406, wire_635, 1'b0, wire_636, NbarT, Si, 1'b0);
dff DFF_77  (wire_75, wire_663, wire_406, wire_661, 1'b0, wire_662, NbarT, Si, 1'b0);
dff DFF_78  (wire_77, wire_664, wire_406, wire_661, 1'b0, wire_662, NbarT, Si, 1'b0);
dff DFF_79  (wire_79, wire_665, wire_406, wire_661, 1'b0, wire_662, NbarT, Si, 1'b0);
dff DFF_80  (wire_81, wire_666, wire_406, wire_661, 1'b0, wire_662, NbarT, Si, 1'b0);
dff DFF_81  (wire_83, wire_667, wire_406, wire_661, 1'b0, wire_662, NbarT, Si, 1'b0);
dff DFF_82  (wire_85, wire_668, wire_406, wire_661, 1'b0, wire_662, NbarT, Si, 1'b0);
dff DFF_83  (wire_87, wire_669, wire_406, wire_661, 1'b0, wire_662, NbarT, Si, 1'b0);
dff DFF_84  (wire_89, wire_670, wire_406, wire_661, 1'b0, wire_662, NbarT, Si, 1'b0);

endmodule
