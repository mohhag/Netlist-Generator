
//Verilog file of module mult8


`timescale 1 ns / 1ns

module mult8_net(i1,
i2,
o);
input [0:7]i1;
input [0:7]i2;
output [0:7]o;
wire
wire_1,
wire_2,
wire_3,
wire_4,
wire_5,
wire_6,
wire_7,
wire_8,
wire_9,
wire_10,
wire_11,
wire_12,
wire_13,
wire_14,
wire_15,
wire_16,
wire_17,
wire_18,
wire_19,
wire_20,
wire_21,
wire_22,
wire_23,
wire_24,
wire_25,
wire_26,
wire_27,
wire_28,
wire_29,
wire_30,
wire_31,
wire_32,
wire_33,
wire_34,
wire_35,
wire_36,
wire_37,
wire_38,
wire_39,
wire_40,
wire_41,
wire_42,
wire_43,
wire_44,
wire_45,
wire_46,
wire_47,
wire_48,
wire_49,
wire_50,
wire_51,
wire_52,
wire_53,
wire_54,
wire_55,
wire_56,
wire_57,
wire_58,
wire_59,
wire_60,
wire_61,
wire_62,
wire_63,
wire_64,
wire_65,
wire_66,
wire_67,
wire_68,
wire_69,
wire_70,
wire_71,
wire_72,
wire_73,
wire_74,
wire_75,
wire_76,
wire_77,
wire_78,
wire_79,
wire_80,
wire_81,
wire_82,
wire_83,
wire_84,
wire_85,
wire_86,
wire_87,
wire_88,
wire_89,
wire_90,
wire_91,
wire_92,
wire_93,
wire_94,
wire_95,
wire_96,
wire_97,
wire_98,
wire_99,
wire_100,
wire_101,
wire_102,
wire_103,
wire_104,
wire_105,
wire_106,
wire_107,
wire_108,
wire_109,
wire_110,
wire_111,
wire_112,
wire_113,
wire_114,
wire_115,
wire_116,
wire_117,
wire_118,
wire_119,
wire_120,
wire_121,
wire_122,
wire_123,
wire_124,
wire_125,
wire_126,
wire_127,
wire_128,
wire_129,
wire_130,
wire_131,
wire_132,
wire_133,
wire_134,
wire_135,
wire_136,
wire_137,
wire_138,
wire_139,
wire_140,
wire_141,
wire_142,
wire_143,
wire_144,
wire_145,
wire_146,
wire_147,
wire_148,
wire_149,
wire_150,
wire_151,
wire_152,
wire_153,
wire_154,
wire_155,
wire_156,
wire_157,
wire_158,
wire_159,
wire_160,
wire_161,
wire_162,
wire_163,
wire_164,
wire_165,
wire_166,
wire_167,
wire_18_0,
wire_18_1,
wire_32_0,
wire_32_1,
wire_32_2,
wire_15_0,
wire_15_1,
wire_40_0,
wire_40_1,
wire_40_2,
wire_44_0,
wire_44_1,
wire_44_2,
wire_12_0,
wire_12_1,
wire_52_0,
wire_52_1,
wire_52_2,
wire_56_0,
wire_56_1,
wire_56_2,
wire_60_0,
wire_60_1,
wire_60_2,
wire_9_0,
wire_9_1,
wire_68_0,
wire_68_1,
wire_68_2,
wire_72_0,
wire_72_1,
wire_72_2,
wire_76_0,
wire_76_1,
wire_76_2,
wire_80_0,
wire_80_1,
wire_80_2,
wire_6_0,
wire_6_1,
wire_79_0,
wire_79_1,
wire_79_2,
wire_59_0,
wire_59_1,
wire_59_2,
wire_43_0,
wire_43_1,
wire_43_2,
wire_31_0,
wire_31_1,
wire_31_2,
wire_88_0,
wire_88_1,
wire_88_2,
wire_92_0,
wire_92_1,
wire_96_0,
wire_96_1,
wire_100_0,
wire_100_1,
wire_104_0,
wire_104_1,
wire_103_0,
wire_103_1,
wire_103_2,
wire_3_0,
wire_3_1,
wire_89_0,
wire_89_1,
wire_89_2,
wire_93_0,
wire_93_1,
wire_93_2,
wire_97_0,
wire_97_1,
wire_97_2,
wire_101_0,
wire_101_1,
wire_101_2,
wire_105_0,
wire_105_1,
wire_105_2,
wire_2_0,
wire_2_1,
wire_69_0,
wire_69_1,
wire_73_0,
wire_73_1,
wire_77_0,
wire_77_1,
wire_81_0,
wire_81_1,
wire_5_0,
wire_5_1,
wire_53_0,
wire_53_1,
wire_57_0,
wire_57_1,
wire_61_0,
wire_61_1,
wire_8_0,
wire_8_1,
wire_41_0,
wire_41_1,
wire_45_0,
wire_45_1,
wire_11_0,
wire_11_1,
wire_33_0,
wire_33_1,
wire_14_0,
wire_14_1,
wire_17_0,
wire_17_1,
wire_99_0,
wire_99_1,
wire_99_2,
wire_95_0,
wire_95_1,
wire_95_2,
wire_91_0,
wire_91_1,
wire_91_2,
wire_87_0,
wire_87_1,
wire_87_2,
wire_75_0,
wire_75_1,
wire_75_2,
wire_71_0,
wire_71_1,
wire_71_2,
wire_67_0,
wire_67_1,
wire_67_2,
wire_55_0,
wire_55_1,
wire_55_2,
wire_51_0,
wire_51_1,
wire_51_2,
wire_39_0,
wire_39_1,
wire_39_2,
wire_150_0,
wire_150_1,
wire_150_2,
wire_150_3,
wire_150_4,
wire_150_5,
wire_150_6,
wire_150_7,
wire_143_0,
wire_143_1,
wire_143_2,
wire_143_3,
wire_143_4,
wire_143_5,
wire_143_6,
wire_140_0,
wire_140_1,
wire_140_2,
wire_140_3,
wire_140_4,
wire_140_5,
wire_137_0,
wire_137_1,
wire_137_2,
wire_137_3,
wire_137_4,
wire_134_0,
wire_134_1,
wire_134_2,
wire_134_3,
wire_131_0,
wire_131_1,
wire_131_2,
wire_130_0,
wire_130_1,
wire_127_0,
wire_127_1,
wire_127_2,
wire_127_3,
wire_127_4,
wire_127_5,
wire_127_6,
wire_127_7,
wire_144_0,
wire_144_1,
wire_144_2,
wire_144_3,
wire_144_4,
wire_144_5,
wire_144_6,
wire_151_0,
wire_151_1,
wire_151_2,
wire_151_3,
wire_151_4,
wire_151_5,
wire_156_0,
wire_156_1,
wire_156_2,
wire_156_3,
wire_156_4,
wire_160_0,
wire_160_1,
wire_160_2,
wire_160_3,
wire_163_0,
wire_163_1,
wire_163_2,
wire_165_0,
wire_165_1;

pin #(16) pin_0 ({i1[0], i1[1], i1[2], i1[3], i1[4], i1[5], i1[6], i1[7], i2[0], i2[1], i2[2], i2[3], i2[4], i2[5], i2[6], i2[7]}, {i1_0, i1_1, i1_2, i1_3, i1_4, i1_5, i1_6, i1_7, i2_0, i2_1, i2_2, i2_3, i2_4, i2_5, i2_6, i2_7});

pout #(8) pout_0 ({o_0, o_1, o_2, o_3, o_4, o_5, o_6, o_7}, {o[0], o[1], o[2], o[3], o[4], o[5], o[6], o[7]});

fanout_n #(2, 0, 0) FANOUT_1 (wire_18, {wire_18_0, wire_18_1});
fanout_n #(3, 0, 0) FANOUT_2 (wire_32, {wire_32_0, wire_32_1, wire_32_2});
fanout_n #(2, 0, 0) FANOUT_3 (wire_15, {wire_15_0, wire_15_1});
fanout_n #(3, 0, 0) FANOUT_4 (wire_40, {wire_40_0, wire_40_1, wire_40_2});
fanout_n #(3, 0, 0) FANOUT_5 (wire_44, {wire_44_0, wire_44_1, wire_44_2});
fanout_n #(2, 0, 0) FANOUT_6 (wire_12, {wire_12_0, wire_12_1});
fanout_n #(3, 0, 0) FANOUT_7 (wire_52, {wire_52_0, wire_52_1, wire_52_2});
fanout_n #(3, 0, 0) FANOUT_8 (wire_56, {wire_56_0, wire_56_1, wire_56_2});
fanout_n #(3, 0, 0) FANOUT_9 (wire_60, {wire_60_0, wire_60_1, wire_60_2});
fanout_n #(2, 0, 0) FANOUT_10 (wire_9, {wire_9_0, wire_9_1});
fanout_n #(3, 0, 0) FANOUT_11 (wire_68, {wire_68_0, wire_68_1, wire_68_2});
fanout_n #(3, 0, 0) FANOUT_12 (wire_72, {wire_72_0, wire_72_1, wire_72_2});
fanout_n #(3, 0, 0) FANOUT_13 (wire_76, {wire_76_0, wire_76_1, wire_76_2});
fanout_n #(3, 0, 0) FANOUT_14 (wire_80, {wire_80_0, wire_80_1, wire_80_2});
fanout_n #(2, 0, 0) FANOUT_15 (wire_6, {wire_6_0, wire_6_1});
fanout_n #(3, 0, 0) FANOUT_16 (wire_79, {wire_79_0, wire_79_1, wire_79_2});
fanout_n #(3, 0, 0) FANOUT_17 (wire_59, {wire_59_0, wire_59_1, wire_59_2});
fanout_n #(3, 0, 0) FANOUT_18 (wire_43, {wire_43_0, wire_43_1, wire_43_2});
fanout_n #(3, 0, 0) FANOUT_19 (wire_31, {wire_31_0, wire_31_1, wire_31_2});
fanout_n #(3, 0, 0) FANOUT_20 (wire_88, {wire_88_0, wire_88_1, wire_88_2});
fanout_n #(2, 0, 0) FANOUT_21 (wire_92, {wire_92_0, wire_92_1});
fanout_n #(2, 0, 0) FANOUT_22 (wire_96, {wire_96_0, wire_96_1});
fanout_n #(2, 0, 0) FANOUT_23 (wire_100, {wire_100_0, wire_100_1});
fanout_n #(2, 0, 0) FANOUT_24 (wire_104, {wire_104_0, wire_104_1});
fanout_n #(3, 0, 0) FANOUT_25 (wire_103, {wire_103_0, wire_103_1, wire_103_2});
fanout_n #(2, 0, 0) FANOUT_26 (wire_3, {wire_3_0, wire_3_1});
fanout_n #(3, 0, 0) FANOUT_27 (wire_89, {wire_89_0, wire_89_1, wire_89_2});
fanout_n #(3, 0, 0) FANOUT_28 (wire_93, {wire_93_0, wire_93_1, wire_93_2});
fanout_n #(3, 0, 0) FANOUT_29 (wire_97, {wire_97_0, wire_97_1, wire_97_2});
fanout_n #(3, 0, 0) FANOUT_30 (wire_101, {wire_101_0, wire_101_1, wire_101_2});
fanout_n #(3, 0, 0) FANOUT_31 (wire_105, {wire_105_0, wire_105_1, wire_105_2});
fanout_n #(2, 0, 0) FANOUT_32 (wire_2, {wire_2_0, wire_2_1});
fanout_n #(2, 0, 0) FANOUT_33 (wire_69, {wire_69_0, wire_69_1});
fanout_n #(2, 0, 0) FANOUT_34 (wire_73, {wire_73_0, wire_73_1});
fanout_n #(2, 0, 0) FANOUT_35 (wire_77, {wire_77_0, wire_77_1});
fanout_n #(2, 0, 0) FANOUT_36 (wire_81, {wire_81_0, wire_81_1});
fanout_n #(2, 0, 0) FANOUT_37 (wire_5, {wire_5_0, wire_5_1});
fanout_n #(2, 0, 0) FANOUT_38 (wire_53, {wire_53_0, wire_53_1});
fanout_n #(2, 0, 0) FANOUT_39 (wire_57, {wire_57_0, wire_57_1});
fanout_n #(2, 0, 0) FANOUT_40 (wire_61, {wire_61_0, wire_61_1});
fanout_n #(2, 0, 0) FANOUT_41 (wire_8, {wire_8_0, wire_8_1});
fanout_n #(2, 0, 0) FANOUT_42 (wire_41, {wire_41_0, wire_41_1});
fanout_n #(2, 0, 0) FANOUT_43 (wire_45, {wire_45_0, wire_45_1});
fanout_n #(2, 0, 0) FANOUT_44 (wire_11, {wire_11_0, wire_11_1});
fanout_n #(2, 0, 0) FANOUT_45 (wire_33, {wire_33_0, wire_33_1});
fanout_n #(2, 0, 0) FANOUT_46 (wire_14, {wire_14_0, wire_14_1});
fanout_n #(2, 0, 0) FANOUT_47 (wire_17, {wire_17_0, wire_17_1});
fanout_n #(3, 0, 0) FANOUT_48 (wire_99, {wire_99_0, wire_99_1, wire_99_2});
fanout_n #(3, 0, 0) FANOUT_49 (wire_95, {wire_95_0, wire_95_1, wire_95_2});
fanout_n #(3, 0, 0) FANOUT_50 (wire_91, {wire_91_0, wire_91_1, wire_91_2});
fanout_n #(3, 0, 0) FANOUT_51 (wire_87, {wire_87_0, wire_87_1, wire_87_2});
fanout_n #(3, 0, 0) FANOUT_52 (wire_75, {wire_75_0, wire_75_1, wire_75_2});
fanout_n #(3, 0, 0) FANOUT_53 (wire_71, {wire_71_0, wire_71_1, wire_71_2});
fanout_n #(3, 0, 0) FANOUT_54 (wire_67, {wire_67_0, wire_67_1, wire_67_2});
fanout_n #(3, 0, 0) FANOUT_55 (wire_55, {wire_55_0, wire_55_1, wire_55_2});
fanout_n #(3, 0, 0) FANOUT_56 (wire_51, {wire_51_0, wire_51_1, wire_51_2});
fanout_n #(3, 0, 0) FANOUT_57 (wire_39, {wire_39_0, wire_39_1, wire_39_2});
fanout_n #(8, 0, 0) FANOUT_58 (wire_150, {wire_150_0, wire_150_1, wire_150_2, wire_150_3, wire_150_4, wire_150_5, wire_150_6, wire_150_7});
fanout_n #(7, 0, 0) FANOUT_59 (wire_143, {wire_143_0, wire_143_1, wire_143_2, wire_143_3, wire_143_4, wire_143_5, wire_143_6});
fanout_n #(6, 0, 0) FANOUT_60 (wire_140, {wire_140_0, wire_140_1, wire_140_2, wire_140_3, wire_140_4, wire_140_5});
fanout_n #(5, 0, 0) FANOUT_61 (wire_137, {wire_137_0, wire_137_1, wire_137_2, wire_137_3, wire_137_4});
fanout_n #(4, 0, 0) FANOUT_62 (wire_134, {wire_134_0, wire_134_1, wire_134_2, wire_134_3});
fanout_n #(3, 0, 0) FANOUT_63 (wire_131, {wire_131_0, wire_131_1, wire_131_2});
fanout_n #(2, 0, 0) FANOUT_64 (wire_130, {wire_130_0, wire_130_1});
fanout_n #(8, 0, 0) FANOUT_65 (wire_127, {wire_127_0, wire_127_1, wire_127_2, wire_127_3, wire_127_4, wire_127_5, wire_127_6, wire_127_7});
fanout_n #(7, 0, 0) FANOUT_66 (wire_144, {wire_144_0, wire_144_1, wire_144_2, wire_144_3, wire_144_4, wire_144_5, wire_144_6});
fanout_n #(6, 0, 0) FANOUT_67 (wire_151, {wire_151_0, wire_151_1, wire_151_2, wire_151_3, wire_151_4, wire_151_5});
fanout_n #(5, 0, 0) FANOUT_68 (wire_156, {wire_156_0, wire_156_1, wire_156_2, wire_156_3, wire_156_4});
fanout_n #(4, 0, 0) FANOUT_69 (wire_160, {wire_160_0, wire_160_1, wire_160_2, wire_160_3});
fanout_n #(3, 0, 0) FANOUT_70 (wire_163, {wire_163_0, wire_163_1, wire_163_2});
fanout_n #(2, 0, 0) FANOUT_71 (wire_165, {wire_165_0, wire_165_1});


xor_n #(2, 0, 0) XOR_1 (wire_1, {wire_2_0, wire_3_0});
xor_n #(2, 0, 0) XOR_2 (wire_4, {wire_5_0, wire_6_0});
xor_n #(2, 0, 0) XOR_3 (wire_7, {wire_8_0, wire_9_0});
xor_n #(2, 0, 0) XOR_4 (wire_10, {wire_11_0, wire_12_0});
xor_n #(2, 0, 0) XOR_5 (wire_13, {wire_14_0, wire_15_0});
xor_n #(2, 0, 0) XOR_6 (wire_16, {wire_17_0, wire_18_0});
xor_n #(2, 0, 0) XOR_7 (wire_19, {wire_20, wire_21});
xor_n #(2, 0, 0) XOR_8 (wire_21, {wire_22, wire_23});
xor_n #(2, 0, 0) XOR_9 (wire_22, {wire_24, wire_25});
xor_n #(2, 0, 0) XOR_10 (wire_24, {wire_26, wire_27});
xor_n #(2, 0, 0) XOR_11 (wire_26, {wire_28, wire_29});
xor_n #(2, 0, 0) XOR_12 (wire_18, {wire_30, wire_31_0});
xor_n #(2, 0, 0) XOR_13 (wire_30, {wire_32_0, wire_33_0});
xor_n #(2, 0, 0) XOR_14 (wire_28, {wire_34, wire_35});
xor_n #(2, 0, 0) XOR_15 (wire_34, {wire_36, wire_37});
xor_n #(2, 0, 0) XOR_16 (wire_32, {wire_38, wire_39_0});
xor_n #(2, 0, 0) XOR_17 (wire_38, {wire_40_0, wire_41_0});
xor_n #(2, 0, 0) XOR_18 (wire_15, {wire_42, wire_43_0});
xor_n #(2, 0, 0) XOR_19 (wire_42, {wire_44_0, wire_45_0});
xor_n #(2, 0, 0) XOR_20 (wire_36, {wire_46, wire_47});
xor_n #(2, 0, 0) XOR_21 (wire_46, {wire_48, wire_49});
xor_n #(2, 0, 0) XOR_22 (wire_40, {wire_50, wire_51_0});
xor_n #(2, 0, 0) XOR_23 (wire_50, {wire_52_0, wire_53_0});
xor_n #(2, 0, 0) XOR_24 (wire_44, {wire_54, wire_55_0});
xor_n #(2, 0, 0) XOR_25 (wire_54, {wire_56_0, wire_57_0});
xor_n #(2, 0, 0) XOR_26 (wire_12, {wire_58, wire_59_0});
xor_n #(2, 0, 0) XOR_27 (wire_58, {wire_60_0, wire_61_0});
xor_n #(2, 0, 0) XOR_28 (wire_48, {wire_62, wire_63});
xor_n #(2, 0, 0) XOR_29 (wire_62, {wire_64, wire_65});
xor_n #(2, 0, 0) XOR_30 (wire_52, {wire_66, wire_67_0});
xor_n #(2, 0, 0) XOR_31 (wire_66, {wire_68_0, wire_69_0});
xor_n #(2, 0, 0) XOR_32 (wire_56, {wire_70, wire_71_0});
xor_n #(2, 0, 0) XOR_33 (wire_70, {wire_72_0, wire_73_0});
xor_n #(2, 0, 0) XOR_34 (wire_60, {wire_74, wire_75_0});
xor_n #(2, 0, 0) XOR_35 (wire_74, {wire_76_0, wire_77_0});
xor_n #(2, 0, 0) XOR_36 (wire_9, {wire_78, wire_79_0});
xor_n #(2, 0, 0) XOR_37 (wire_78, {wire_80_0, wire_81_0});
xor_n #(2, 0, 0) XOR_38 (wire_64, {wire_82, wire_83});
xor_n #(2, 0, 0) XOR_39 (wire_82, {wire_84, wire_85});
xor_n #(2, 0, 0) XOR_40 (wire_68, {wire_86, wire_87_0});
xor_n #(2, 0, 0) XOR_41 (wire_86, {wire_88_0, wire_89_0});
xor_n #(2, 0, 0) XOR_42 (wire_72, {wire_90, wire_91_0});
xor_n #(2, 0, 0) XOR_43 (wire_90, {wire_92_0, wire_93_0});
xor_n #(2, 0, 0) XOR_44 (wire_76, {wire_94, wire_95_0});
xor_n #(2, 0, 0) XOR_45 (wire_94, {wire_96_0, wire_97_0});
xor_n #(2, 0, 0) XOR_46 (wire_80, {wire_98, wire_99_0});
xor_n #(2, 0, 0) XOR_47 (wire_98, {wire_100_0, wire_101_0});
xor_n #(2, 0, 0) XOR_48 (wire_6, {wire_102, wire_103_0});
xor_n #(2, 0, 0) XOR_49 (wire_102, {wire_104_0, wire_105_0});
and_n #(2, 0, 0) AND_1 (wire_79, {wire_6_1, wire_5_1});
and_n #(2, 0, 0) AND_2 (wire_106, {wire_80_1, wire_79_1});
or_n #(2, 0, 0) OR_1 (wire_107, {wire_80_2, wire_79_2});
and_n #(2, 0, 0) AND_3 (wire_108, {wire_76_1, wire_75_1});
or_n #(2, 0, 0) OR_2 (wire_109, {wire_76_2, wire_75_2});
and_n #(2, 0, 0) AND_4 (wire_110, {wire_72_1, wire_71_1});
or_n #(2, 0, 0) OR_3 (wire_111, {wire_72_2, wire_71_2});
and_n #(2, 0, 0) AND_5 (wire_112, {wire_68_1, wire_67_1});
or_n #(2, 0, 0) OR_4 (wire_113, {wire_68_2, wire_67_2});
and_n #(2, 0, 0) AND_6 (wire_59, {wire_9_1, wire_8_1});
and_n #(2, 0, 0) AND_7 (wire_114, {wire_60_1, wire_59_1});
or_n #(2, 0, 0) OR_5 (wire_115, {wire_60_2, wire_59_2});
and_n #(2, 0, 0) AND_8 (wire_116, {wire_56_1, wire_55_1});
or_n #(2, 0, 0) OR_6 (wire_117, {wire_56_2, wire_55_2});
and_n #(2, 0, 0) AND_9 (wire_118, {wire_52_1, wire_51_1});
or_n #(2, 0, 0) OR_7 (wire_119, {wire_52_2, wire_51_2});
and_n #(2, 0, 0) AND_10 (wire_43, {wire_12_1, wire_11_1});
and_n #(2, 0, 0) AND_11 (wire_120, {wire_44_1, wire_43_1});
or_n #(2, 0, 0) OR_8 (wire_121, {wire_44_2, wire_43_2});
and_n #(2, 0, 0) AND_12 (wire_122, {wire_40_1, wire_39_1});
or_n #(2, 0, 0) OR_9 (wire_123, {wire_40_2, wire_39_2});
and_n #(2, 0, 0) AND_13 (wire_31, {wire_15_1, wire_14_1});
and_n #(2, 0, 0) AND_14 (wire_124, {wire_32_1, wire_31_1});
or_n #(2, 0, 0) OR_10 (wire_125, {wire_32_2, wire_31_2});
and_n #(2, 0, 0) AND_15 (wire_23, {wire_18_1, wire_17_1});
and_n #(2, 0, 0) AND_16 (wire_84, {wire_126, wire_127_0});
and_n #(2, 0, 0) AND_17 (wire_128, {wire_88_1, wire_87_1});
and_n #(2, 0, 0) AND_18 (wire_129, {wire_88_2, wire_89_1});
and_n #(2, 0, 0) AND_19 (wire_88, {wire_130_0, wire_127_1});
and_n #(2, 0, 0) AND_20 (wire_92, {wire_131_0, wire_127_2});
and_n #(2, 0, 0) AND_21 (wire_132, {wire_92_1, wire_133});
and_n #(2, 0, 0) AND_22 (wire_96, {wire_134_0, wire_127_3});
and_n #(2, 0, 0) AND_23 (wire_135, {wire_96_1, wire_136});
and_n #(2, 0, 0) AND_24 (wire_100, {wire_137_0, wire_127_4});
and_n #(2, 0, 0) AND_25 (wire_138, {wire_100_1, wire_139});
and_n #(2, 0, 0) AND_26 (wire_104, {wire_140_0, wire_127_5});
and_n #(2, 0, 0) AND_27 (wire_141, {wire_104_1, wire_142});
and_n #(2, 0, 0) AND_28 (wire_103, {wire_3_1, wire_2_1});
and_n #(2, 0, 0) AND_29 (wire_3, {wire_143_0, wire_127_6});
and_n #(2, 0, 0) AND_30 (wire_85, {wire_130_1, wire_144_0});
and_n #(2, 0, 0) AND_31 (wire_145, {wire_89_2, wire_87_2});
and_n #(2, 0, 0) AND_32 (wire_89, {wire_131_1, wire_144_1});
and_n #(2, 0, 0) AND_33 (wire_93, {wire_134_1, wire_144_2});
and_n #(2, 0, 0) AND_34 (wire_146, {wire_93_1, wire_91_1});
or_n #(2, 0, 0) OR_11 (wire_133, {wire_93_2, wire_91_2});
and_n #(2, 0, 0) AND_35 (wire_97, {wire_137_1, wire_144_3});
and_n #(2, 0, 0) AND_36 (wire_147, {wire_97_1, wire_95_1});
or_n #(2, 0, 0) OR_12 (wire_136, {wire_97_2, wire_95_2});
and_n #(2, 0, 0) AND_37 (wire_101, {wire_140_1, wire_144_4});
and_n #(2, 0, 0) AND_38 (wire_148, {wire_101_1, wire_99_1});
or_n #(2, 0, 0) OR_13 (wire_139, {wire_101_2, wire_99_2});
and_n #(2, 0, 0) AND_39 (wire_105, {wire_143_1, wire_144_5});
and_n #(2, 0, 0) AND_40 (wire_149, {wire_105_1, wire_103_1});
or_n #(2, 0, 0) OR_14 (wire_142, {wire_105_2, wire_103_2});
and_n #(2, 0, 0) AND_41 (wire_2, {wire_150_0, wire_144_6});
and_n #(2, 0, 0) AND_42 (wire_65, {wire_131_2, wire_151_0});
and_n #(2, 0, 0) AND_43 (wire_69, {wire_134_2, wire_151_1});
and_n #(2, 0, 0) AND_44 (wire_152, {wire_69_1, wire_113});
and_n #(2, 0, 0) AND_45 (wire_73, {wire_137_2, wire_151_2});
and_n #(2, 0, 0) AND_46 (wire_153, {wire_73_1, wire_111});
and_n #(2, 0, 0) AND_47 (wire_77, {wire_140_2, wire_151_3});
and_n #(2, 0, 0) AND_48 (wire_154, {wire_77_1, wire_109});
and_n #(2, 0, 0) AND_49 (wire_81, {wire_143_2, wire_151_4});
and_n #(2, 0, 0) AND_50 (wire_155, {wire_81_1, wire_107});
and_n #(2, 0, 0) AND_51 (wire_5, {wire_150_1, wire_151_5});
and_n #(2, 0, 0) AND_52 (wire_49, {wire_134_3, wire_156_0});
and_n #(2, 0, 0) AND_53 (wire_53, {wire_137_3, wire_156_1});
and_n #(2, 0, 0) AND_54 (wire_157, {wire_53_1, wire_119});
and_n #(2, 0, 0) AND_55 (wire_57, {wire_140_3, wire_156_2});
and_n #(2, 0, 0) AND_56 (wire_158, {wire_57_1, wire_117});
and_n #(2, 0, 0) AND_57 (wire_61, {wire_143_3, wire_156_3});
and_n #(2, 0, 0) AND_58 (wire_159, {wire_61_1, wire_115});
and_n #(2, 0, 0) AND_59 (wire_8, {wire_150_2, wire_156_4});
and_n #(2, 0, 0) AND_60 (wire_37, {wire_137_4, wire_160_0});
and_n #(2, 0, 0) AND_61 (wire_41, {wire_140_4, wire_160_1});
and_n #(2, 0, 0) AND_62 (wire_161, {wire_41_1, wire_123});
and_n #(2, 0, 0) AND_63 (wire_45, {wire_143_4, wire_160_2});
and_n #(2, 0, 0) AND_64 (wire_162, {wire_45_1, wire_121});
and_n #(2, 0, 0) AND_65 (wire_11, {wire_150_3, wire_160_3});
and_n #(2, 0, 0) AND_66 (wire_29, {wire_140_5, wire_163_0});
and_n #(2, 0, 0) AND_67 (wire_33, {wire_143_5, wire_163_1});
and_n #(2, 0, 0) AND_68 (wire_164, {wire_33_1, wire_125});
and_n #(2, 0, 0) AND_69 (wire_14, {wire_150_4, wire_163_2});
and_n #(2, 0, 0) AND_70 (wire_25, {wire_143_6, wire_165_0});
and_n #(2, 0, 0) AND_71 (wire_17, {wire_150_5, wire_165_1});
and_n #(2, 0, 0) AND_72 (wire_20, {wire_150_6, wire_166});
or_n #(2, 0, 0) OR_15 (wire_99, {wire_149, wire_141});
or_n #(2, 0, 0) OR_16 (wire_95, {wire_148, wire_138});
or_n #(2, 0, 0) OR_17 (wire_91, {wire_147, wire_135});
or_n #(2, 0, 0) OR_18 (wire_87, {wire_146, wire_132});
or_n #(3, 0, 0) OR_19 (wire_83, {wire_129, wire_128, wire_145});
or_n #(2, 0, 0) OR_20 (wire_75, {wire_106, wire_155});
or_n #(2, 0, 0) OR_21 (wire_71, {wire_108, wire_154});
or_n #(2, 0, 0) OR_22 (wire_67, {wire_110, wire_153});
or_n #(2, 0, 0) OR_23 (wire_63, {wire_112, wire_152});
or_n #(2, 0, 0) OR_24 (wire_55, {wire_114, wire_159});
or_n #(2, 0, 0) OR_25 (wire_51, {wire_116, wire_158});
or_n #(2, 0, 0) OR_26 (wire_47, {wire_118, wire_157});
or_n #(2, 0, 0) OR_27 (wire_39, {wire_120, wire_162});
or_n #(2, 0, 0) OR_28 (wire_35, {wire_122, wire_161});
or_n #(2, 0, 0) OR_29 (wire_27, {wire_124, wire_164});
bufg #(0, 0) BUF_1 (wire_150, i1_7);
bufg #(0, 0) BUF_2 (wire_143, i1_6);
bufg #(0, 0) BUF_3 (wire_140, i1_5);
bufg #(0, 0) BUF_4 (wire_137, i1_4);
bufg #(0, 0) BUF_5 (wire_134, i1_3);
bufg #(0, 0) BUF_6 (wire_131, i1_2);
bufg #(0, 0) BUF_7 (wire_130, i1_1);
bufg #(0, 0) BUF_8 (wire_126, i1_0);
and_n #(2, 0, 0) AND_73 (wire_167, {wire_150_7, wire_127_7});
bufg #(0, 0) BUF_9 (wire_127, i2_7);
bufg #(0, 0) BUF_10 (wire_144, i2_6);
bufg #(0, 0) BUF_11 (wire_151, i2_5);
bufg #(0, 0) BUF_12 (wire_156, i2_4);
bufg #(0, 0) BUF_13 (wire_160, i2_3);
bufg #(0, 0) BUF_14 (wire_163, i2_2);
bufg #(0, 0) BUF_15 (wire_165, i2_1);
bufg #(0, 0) BUF_16 (wire_166, i2_0);
bufg #(0, 0) BUF_17 (o_7, wire_167);
bufg #(0, 0) BUF_18 (o_6, wire_1);
bufg #(0, 0) BUF_19 (o_5, wire_4);
bufg #(0, 0) BUF_20 (o_4, wire_7);
bufg #(0, 0) BUF_21 (o_3, wire_10);
bufg #(0, 0) BUF_22 (o_2, wire_13);
bufg #(0, 0) BUF_23 (o_1, wire_16);
bufg #(0, 0) BUF_24 (o_0, wire_19);

endmodule
